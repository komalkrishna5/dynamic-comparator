magic
tech sky130A
magscale 1 2
timestamp 1646259600
<< error_p >>
rect -159 222 -129 226
rect -63 222 -33 226
rect 33 222 63 226
rect 129 222 159 226
rect -217 144 -159 200
rect -221 -144 -159 144
rect -217 -200 -159 -144
rect -129 -200 -63 200
rect -33 -200 33 200
rect 63 -200 129 200
rect 159 144 217 200
rect 159 -144 221 144
rect 159 -200 217 -144
rect -159 -226 -129 -222
rect -63 -226 -33 -222
rect 33 -226 63 -222
rect 129 -226 159 -222
<< nmos >>
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
<< ndiff >>
rect -217 144 -159 200
rect -221 132 -159 144
rect -221 -132 -209 132
rect -175 -132 -159 132
rect -221 -144 -159 -132
rect -217 -200 -159 -144
rect -129 132 -63 200
rect -129 -132 -113 132
rect -79 -132 -63 132
rect -129 -200 -63 -132
rect -33 132 33 200
rect -33 -132 -17 132
rect 17 -132 33 132
rect -33 -200 33 -132
rect 63 132 129 200
rect 63 -132 79 132
rect 113 -132 129 132
rect 63 -200 129 -132
rect 159 144 217 200
rect 159 132 221 144
rect 159 -132 175 132
rect 209 -132 221 132
rect 159 -144 221 -132
rect 159 -200 217 -144
<< ndiffc >>
rect -209 -132 -175 132
rect -113 -132 -79 132
rect -17 -132 17 132
rect 79 -132 113 132
rect 175 -132 209 132
<< poly >>
rect -159 200 -129 222
rect -63 200 -33 222
rect 33 200 63 222
rect 129 200 159 222
rect -159 -222 -129 -200
rect -63 -222 -33 -200
rect 33 -222 63 -200
rect 129 -222 159 -200
<< locali >>
rect -209 132 -175 148
rect -209 -148 -175 -132
rect -113 132 -79 148
rect -113 -148 -79 -132
rect -17 132 17 148
rect -17 -148 17 -132
rect 79 132 113 148
rect 79 -148 113 -132
rect 175 132 209 148
rect 175 -148 209 -132
<< viali >>
rect -209 -132 -175 132
rect -113 -132 -79 132
rect -17 -132 17 132
rect 79 -132 113 132
rect 175 -132 209 132
<< metal1 >>
rect -215 132 -169 144
rect -215 -132 -209 132
rect -175 -132 -169 132
rect -215 -144 -169 -132
rect -119 132 -73 144
rect -119 -132 -113 132
rect -79 -132 -73 132
rect -119 -144 -73 -132
rect -23 132 23 144
rect -23 -132 -17 132
rect 17 -132 23 132
rect -23 -144 23 -132
rect 73 132 119 144
rect 73 -132 79 132
rect 113 -132 119 132
rect 73 -144 119 -132
rect 169 132 215 144
rect 169 -132 175 132
rect 209 -132 215 132
rect 169 -144 215 -132
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 4 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
