magic
tech sky130A
magscale 1 2
timestamp 1646429429
<< nmos >>
rect -63 -100 -33 100
rect 33 -100 63 100
<< ndiff >>
rect -121 74 -63 100
rect -125 62 -63 74
rect -125 -62 -113 62
rect -79 -62 -63 62
rect -125 -74 -63 -62
rect -121 -100 -63 -74
rect -33 62 33 100
rect -33 -62 -17 62
rect 17 -62 33 62
rect -33 -100 33 -62
rect 63 74 121 100
rect 63 62 125 74
rect 63 -62 79 62
rect 113 -62 125 62
rect 63 -74 125 -62
rect 63 -100 121 -74
<< ndiffc >>
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
<< poly >>
rect -63 122 63 154
rect -63 100 -33 122
rect 33 100 63 122
rect -63 -118 -33 -100
rect 33 -118 63 -100
rect -63 -152 63 -118
<< locali >>
rect -113 62 -79 78
rect -113 -78 -79 -62
rect -17 62 17 78
rect -17 -78 17 -62
rect 79 62 113 78
rect 79 -78 113 -62
<< viali >>
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
<< metal1 >>
rect -119 62 -73 74
rect -119 -62 -113 62
rect -79 -62 -73 62
rect -119 -74 -73 -62
rect -23 62 23 74
rect -23 -62 -17 62
rect 17 -62 23 62
rect -23 -74 23 -62
rect 73 62 119 74
rect 73 -62 79 62
rect 113 -62 119 62
rect 73 -74 119 -62
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 2 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
