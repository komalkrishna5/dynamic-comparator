magic
tech sky130A
timestamp 1647352381
<< nwell >>
rect 391 2526 470 2668
rect -174 1576 74 1784
rect 89 1039 812 1201
rect 88 389 203 522
<< psubdiff >>
rect 43 64 79 76
rect 43 -12 79 0
<< nsubdiff >>
rect 405 2635 444 2647
rect 405 2533 444 2545
rect -21 1712 13 1724
rect -21 1638 13 1650
rect 166 1154 208 1166
rect 166 1069 208 1081
rect 97 504 156 516
rect 97 392 156 404
<< psubdiffcont >>
rect 43 0 79 64
<< nsubdiffcont >>
rect 405 2545 444 2635
rect -21 1650 13 1712
rect 166 1081 208 1154
rect 97 404 156 504
<< poly >>
rect 326 2406 341 2410
rect 183 2303 222 2315
rect 183 2279 192 2303
rect 213 2289 222 2303
rect 684 2290 721 2300
rect 684 2289 692 2290
rect 213 2279 341 2289
rect 183 2266 341 2279
rect 524 2266 692 2289
rect 713 2266 721 2290
rect 684 2259 721 2266
rect 380 1934 492 1945
rect 380 1899 414 1934
rect 464 1899 492 1934
rect 380 1739 492 1899
rect 255 1278 292 1288
rect 255 1259 265 1278
rect 283 1259 292 1278
rect 255 1247 292 1259
rect 545 1278 582 1288
rect 545 1259 555 1278
rect 573 1259 582 1278
rect 545 1247 582 1259
rect 265 1174 280 1247
rect 556 1175 571 1247
rect 409 745 424 803
rect 408 661 424 745
rect 407 638 425 661
rect 401 630 435 638
rect 401 609 409 630
rect 429 609 435 630
rect 401 600 435 609
<< polycont >>
rect 192 2279 213 2303
rect 692 2266 713 2290
rect 414 1899 464 1934
rect 265 1259 283 1278
rect 555 1259 573 1278
rect 409 609 429 630
<< locali >>
rect -1296 2676 -675 2757
rect 1668 2727 2266 2778
rect 1668 2707 1714 2727
rect 1667 2705 1714 2707
rect 1306 2704 1714 2705
rect 198 2699 1714 2704
rect -1296 2319 -673 2676
rect 411 2643 440 2687
rect 574 2676 1714 2699
rect 405 2635 444 2643
rect 405 2537 444 2545
rect 1668 2607 1714 2676
rect 1826 2607 2114 2727
rect 2226 2607 2266 2727
rect 257 2426 388 2460
rect 545 2431 595 2468
rect -1296 2146 -1256 2319
rect -1131 2146 -856 2319
rect -731 2254 -673 2319
rect 184 2303 221 2313
rect 184 2279 192 2303
rect 213 2279 221 2303
rect 184 2272 221 2279
rect 684 2290 721 2300
rect 684 2266 692 2290
rect 713 2266 721 2290
rect 684 2259 721 2266
rect -731 2227 212 2254
rect -731 2146 -673 2227
rect -1296 2045 -673 2146
rect -1296 1948 -681 2045
rect -1296 1413 -673 1948
rect 399 1934 477 1946
rect 399 1899 414 1934
rect 464 1899 477 1934
rect 399 1889 477 1899
rect -25 1849 16 1855
rect -25 1819 -19 1849
rect 10 1819 16 1849
rect -25 1811 16 1819
rect 1668 1848 2266 2607
rect -14 1720 5 1811
rect 1668 1728 1714 1848
rect 1826 1728 2114 1848
rect 2226 1728 2266 1848
rect -21 1712 13 1720
rect -21 1642 13 1650
rect 823 1514 851 1564
rect 823 1497 828 1514
rect 846 1497 851 1514
rect 823 1496 851 1497
rect 1159 1424 1335 1449
rect 1159 1422 1193 1424
rect -1296 1240 -1256 1413
rect -1131 1240 -856 1413
rect -731 1382 -673 1413
rect 1160 1386 1193 1422
rect -731 1381 -17 1382
rect -731 1355 42 1381
rect 1159 1358 1193 1386
rect -731 1240 -673 1355
rect -16 1344 42 1355
rect -16 1318 73 1344
rect -16 1317 42 1318
rect -441 1270 -265 1295
rect 1160 1293 1193 1358
rect 1306 1386 1335 1424
rect 1306 1358 1337 1386
rect 1306 1293 1335 1358
rect -441 1268 -407 1270
rect -1296 863 -673 1240
rect -440 1139 -407 1268
rect -294 1139 -265 1270
rect 256 1278 291 1286
rect 256 1259 265 1278
rect 283 1259 291 1278
rect 256 1251 291 1259
rect 546 1278 581 1286
rect 546 1259 555 1278
rect 573 1259 581 1278
rect 1160 1268 1335 1293
rect 1668 1268 2266 1728
rect 546 1251 581 1259
rect 1668 1232 1714 1268
rect 40 1205 140 1232
rect 691 1231 1029 1232
rect 1641 1231 1714 1232
rect 691 1204 1714 1231
rect 1049 1203 1638 1204
rect -440 1114 -265 1139
rect 166 1154 259 1167
rect 208 1081 259 1154
rect 166 1068 259 1081
rect 1668 1148 1714 1204
rect 1826 1148 2114 1268
rect 2226 1148 2266 1268
rect -1296 690 -1256 863
rect -1131 690 -856 863
rect -731 786 -673 863
rect -731 757 166 786
rect 1160 775 1335 800
rect -731 690 -673 757
rect -1296 213 -673 690
rect -440 679 -265 704
rect -440 548 -407 679
rect -294 548 -265 679
rect 1160 666 1193 775
rect 1159 644 1193 666
rect 1306 644 1335 775
rect 401 630 435 638
rect 1159 637 1335 644
rect 401 609 409 630
rect 429 609 435 630
rect 1160 619 1335 637
rect 401 600 435 609
rect 1668 618 2266 1148
rect 1668 570 1714 618
rect 825 569 1159 570
rect 1335 569 1714 570
rect -440 523 -265 548
rect -135 542 31 567
rect 825 541 1714 569
rect 97 504 213 512
rect 156 415 213 504
rect 1668 498 1714 541
rect 1826 498 2114 618
rect 2226 498 2266 618
rect 97 396 156 404
rect -1296 40 -1256 213
rect -1131 40 -856 213
rect -731 119 -673 213
rect -731 93 13 119
rect 60 101 79 115
rect -731 40 -673 93
rect -1296 -442 -673 40
rect 43 64 79 101
rect 43 -8 79 0
rect -440 -51 -265 -26
rect -440 -182 -407 -51
rect -294 -75 -265 -51
rect -294 -182 -265 -161
rect -440 -208 -265 -182
rect 1668 -403 2266 498
rect 1668 -437 2251 -403
<< viali >>
rect 1714 2607 1826 2727
rect 2114 2607 2226 2727
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect 192 2279 213 2303
rect 692 2266 713 2290
rect 414 1899 464 1934
rect -19 1819 10 1849
rect 1714 1728 1826 1848
rect 2114 1728 2226 1848
rect 153 1539 178 1562
rect 692 1539 717 1562
rect 828 1497 846 1514
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect 1193 1293 1306 1424
rect -407 1139 -294 1270
rect 265 1259 283 1278
rect 555 1259 573 1278
rect 1714 1148 1826 1268
rect 2114 1148 2226 1268
rect -1256 690 -1131 863
rect -856 690 -731 863
rect -407 548 -294 679
rect 1193 644 1306 775
rect 409 609 429 630
rect 1714 498 1826 618
rect 2114 498 2226 618
rect -1256 40 -1131 213
rect -856 40 -731 213
rect -407 -182 -294 -51
<< metal1 >>
rect 1679 2727 1857 2757
rect 1679 2607 1714 2727
rect 1826 2607 1857 2727
rect 1679 2574 1857 2607
rect 2078 2727 2257 2757
rect 2078 2607 2114 2727
rect 2226 2607 2257 2727
rect 2078 2574 2257 2607
rect -1285 2319 -1102 2342
rect -1285 2146 -1256 2319
rect -1131 2146 -1102 2319
rect -1285 2113 -1102 2146
rect -885 2319 -702 2342
rect -885 2146 -856 2319
rect -731 2146 -702 2319
rect 184 2305 221 2313
rect -885 2113 -702 2146
rect -105 2303 221 2305
rect -105 2279 192 2303
rect 213 2279 221 2303
rect -105 2277 221 2279
rect -105 1896 -64 2277
rect 184 2272 221 2277
rect 684 2290 721 2300
rect 684 2266 692 2290
rect 713 2267 986 2290
rect 713 2266 721 2267
rect 943 2266 986 2267
rect 684 2259 721 2266
rect 945 1961 986 2266
rect -104 1564 -64 1896
rect 399 1934 477 1946
rect 399 1899 414 1934
rect 464 1899 477 1934
rect 399 1889 477 1899
rect -25 1849 16 1855
rect 402 1851 521 1864
rect 402 1849 433 1851
rect -25 1819 -19 1849
rect 10 1819 433 1849
rect -25 1818 433 1819
rect -25 1811 16 1818
rect 402 1811 433 1818
rect 485 1811 521 1851
rect 402 1800 521 1811
rect 136 1564 187 1572
rect -104 1562 187 1564
rect -104 1539 153 1562
rect 178 1539 187 1562
rect -104 1536 187 1539
rect -1285 1413 -1102 1438
rect -1285 1240 -1256 1413
rect -1131 1240 -1102 1413
rect -1285 1207 -1102 1240
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect -441 1270 -265 1295
rect -441 1139 -407 1270
rect -294 1139 -265 1270
rect -441 1114 -265 1139
rect -1285 863 -1102 888
rect -1285 690 -1256 863
rect -1131 690 -1102 863
rect -1285 657 -1102 690
rect -885 863 -702 888
rect -885 690 -856 863
rect -731 690 -702 863
rect -885 657 -702 690
rect -441 679 -265 704
rect -441 548 -407 679
rect -294 548 -265 679
rect -441 523 -265 548
rect -1285 213 -1102 238
rect -1285 40 -1256 213
rect -1131 40 -1102 213
rect -1285 7 -1102 40
rect -885 213 -702 238
rect -885 40 -856 213
rect -731 40 -702 213
rect -104 199 -64 1536
rect 136 1515 187 1536
rect 684 1562 726 1572
rect 684 1539 692 1562
rect 717 1561 726 1562
rect 946 1561 986 1961
rect 1678 1848 1857 1878
rect 1678 1728 1714 1848
rect 1826 1728 1857 1848
rect 1678 1695 1857 1728
rect 2078 1848 2257 1878
rect 2078 1728 2114 1848
rect 2226 1728 2257 1848
rect 2078 1695 2257 1728
rect 717 1539 987 1561
rect 684 1536 987 1539
rect 684 1530 726 1536
rect 823 1515 852 1520
rect 136 1514 852 1515
rect 136 1497 828 1514
rect 846 1497 852 1514
rect 946 1501 987 1536
rect 136 1496 852 1497
rect 823 1490 852 1496
rect 256 1282 291 1286
rect 256 1256 262 1282
rect 288 1256 291 1282
rect 256 1251 291 1256
rect 546 1282 581 1286
rect 546 1256 552 1282
rect 578 1256 581 1282
rect 546 1251 581 1256
rect -29 965 153 996
rect 601 969 903 1000
rect -29 293 -1 965
rect 130 950 153 965
rect 130 944 152 950
rect 401 634 435 638
rect 401 605 405 634
rect 433 605 435 634
rect 401 600 435 605
rect 875 293 903 969
rect -29 272 20 293
rect 858 272 903 293
rect 947 206 987 1501
rect 1159 1424 1335 1449
rect 1159 1293 1193 1424
rect 1306 1293 1335 1424
rect 1159 1268 1335 1293
rect 1678 1268 1857 1298
rect 1678 1148 1714 1268
rect 1826 1148 1857 1268
rect 1678 1115 1857 1148
rect 2078 1268 2257 1298
rect 2078 1148 2114 1268
rect 2226 1148 2257 1268
rect 2078 1115 2257 1148
rect 1159 775 1335 800
rect 1159 644 1193 775
rect 1306 644 1335 775
rect 1159 619 1335 644
rect 1678 618 1857 649
rect 1678 498 1714 618
rect 1826 498 1857 618
rect 1678 465 1857 498
rect 2078 618 2257 649
rect 2078 498 2114 618
rect 2226 498 2257 618
rect 2078 465 2257 498
rect -104 171 35 199
rect 819 178 987 206
rect -885 7 -702 40
rect -441 -51 -265 -26
rect -441 -182 -407 -51
rect -294 -182 -265 -51
rect 148 -58 295 54
rect 558 -58 708 56
rect -441 -208 -265 -182
<< via1 >>
rect 1714 2607 1826 2727
rect 2114 2607 2226 2727
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect 433 1811 485 1851
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect -407 1139 -294 1270
rect -1256 690 -1131 863
rect -856 690 -731 863
rect -407 548 -294 679
rect -1256 40 -1131 213
rect -856 40 -731 213
rect 1714 1728 1826 1848
rect 2114 1728 2226 1848
rect 262 1278 288 1282
rect 262 1259 265 1278
rect 265 1259 283 1278
rect 283 1259 288 1278
rect 262 1256 288 1259
rect 552 1278 578 1282
rect 552 1259 555 1278
rect 555 1259 573 1278
rect 573 1259 578 1278
rect 552 1256 578 1259
rect 212 603 240 634
rect 405 630 433 634
rect 405 609 409 630
rect 409 609 429 630
rect 429 609 433 630
rect 405 605 433 609
rect 617 605 645 634
rect 1193 1293 1306 1424
rect 1714 1148 1826 1268
rect 2114 1148 2226 1268
rect 1193 659 1306 775
rect 1193 644 1305 659
rect 1714 498 1826 618
rect 2114 498 2226 618
rect -407 -182 -294 -51
rect 406 5 455 49
<< metal2 >>
rect 1664 2727 2266 2778
rect 1664 2607 1714 2727
rect 1826 2607 2114 2727
rect 2226 2607 2266 2727
rect -1285 2319 -1102 2342
rect -1285 2146 -1256 2319
rect -1131 2146 -1102 2319
rect -1285 2113 -1102 2146
rect -885 2319 -702 2342
rect -885 2146 -856 2319
rect -731 2146 -702 2319
rect -885 2113 -702 2146
rect 402 1851 516 1859
rect 402 1811 433 1851
rect 485 1843 516 1851
rect 1664 1848 2266 2607
rect 1664 1843 1714 1848
rect 485 1811 1714 1843
rect 402 1810 1714 1811
rect 402 1801 516 1810
rect 1664 1728 1714 1810
rect 1826 1728 2114 1848
rect 2226 1728 2266 1848
rect -1285 1413 -1102 1438
rect -1285 1240 -1256 1413
rect -1131 1240 -1102 1413
rect -1285 1207 -1102 1240
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect -460 1279 -259 1471
rect 1139 1424 1340 1472
rect 1139 1293 1193 1424
rect 1306 1293 1340 1424
rect 1139 1290 1340 1293
rect 578 1289 1340 1290
rect 255 1282 292 1288
rect 255 1279 262 1282
rect -460 1270 262 1279
rect -460 1139 -407 1270
rect -294 1256 262 1270
rect 288 1256 292 1282
rect -294 1255 292 1256
rect -294 1139 -259 1255
rect 255 1247 292 1255
rect 545 1282 1340 1289
rect 545 1256 552 1282
rect 578 1263 1340 1282
rect 578 1256 582 1263
rect 545 1247 582 1256
rect -460 1046 -259 1139
rect 1139 1048 1340 1263
rect -460 1013 185 1046
rect -1285 863 -1102 888
rect -1285 690 -1256 863
rect -1131 690 -1102 863
rect -1285 657 -1102 690
rect -885 863 -702 888
rect -885 690 -856 863
rect -731 690 -702 863
rect -885 657 -702 690
rect -460 679 -259 1013
rect 660 1012 1340 1048
rect 1139 775 1340 1012
rect 1139 685 1193 775
rect -460 548 -407 679
rect -294 676 -259 679
rect 400 677 436 678
rect 206 676 436 677
rect -294 652 436 676
rect -294 548 -259 652
rect 206 634 243 652
rect 206 603 212 634
rect 240 603 243 634
rect 206 600 243 603
rect 400 634 436 652
rect 617 660 1193 685
rect 617 638 647 660
rect 400 605 405 634
rect 433 605 436 634
rect 400 600 436 605
rect 613 634 647 638
rect 613 605 617 634
rect 645 605 647 634
rect 613 600 647 605
rect 1139 644 1193 660
rect 1306 659 1340 775
rect 1305 644 1340 659
rect -1285 213 -1102 238
rect -1285 40 -1256 213
rect -1131 40 -1102 213
rect -1285 7 -1102 40
rect -885 213 -702 238
rect -885 40 -856 213
rect -731 40 -702 213
rect -885 7 -702 40
rect -460 -51 -259 548
rect -460 -182 -407 -51
rect -294 -105 -259 -51
rect 397 49 464 55
rect 397 5 406 49
rect 455 5 464 49
rect 397 -105 464 5
rect -294 -150 465 -105
rect -294 -182 -259 -150
rect -460 -268 -259 -182
rect 1139 -268 1340 644
rect 1664 1268 2266 1728
rect 1664 1148 1714 1268
rect 1826 1148 2114 1268
rect 2226 1148 2266 1268
rect 1664 618 2266 1148
rect 1664 498 1714 618
rect 1826 498 2114 618
rect 2226 498 2266 618
rect -460 -412 1341 -268
rect 1664 -403 2266 498
rect 1664 -437 2251 -403
<< via2 >>
rect 1714 2607 1826 2727
rect 2114 2607 2226 2727
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect 1714 1728 1826 1848
rect 2114 1728 2226 1848
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect 1193 1293 1306 1424
rect -407 1139 -294 1270
rect -1256 690 -1131 863
rect -856 690 -731 863
rect -407 548 -294 679
rect 1193 659 1306 775
rect 1193 644 1305 659
rect -1256 40 -1131 213
rect -856 40 -731 213
rect -407 -182 -294 -51
rect 1714 1148 1826 1268
rect 2114 1148 2226 1268
rect 1714 498 1826 618
rect 2114 498 2226 618
<< metal3 >>
rect 1679 2727 1857 2757
rect 1679 2607 1714 2727
rect 1826 2607 1857 2727
rect 1679 2574 1857 2607
rect 2078 2727 2257 2757
rect 2078 2607 2114 2727
rect 2226 2607 2257 2727
rect 2078 2574 2257 2607
rect -1285 2319 -1102 2342
rect -1285 2146 -1256 2319
rect -1131 2146 -1102 2319
rect -1285 2113 -1102 2146
rect -885 2319 -702 2342
rect -885 2146 -856 2319
rect -731 2146 -702 2319
rect -885 2113 -702 2146
rect 1678 1848 1857 1878
rect 1678 1728 1714 1848
rect 1826 1728 1857 1848
rect 1678 1695 1857 1728
rect 2078 1848 2257 1878
rect 2078 1728 2114 1848
rect 2226 1728 2257 1848
rect 2078 1695 2257 1728
rect -1285 1413 -1102 1438
rect -1285 1240 -1256 1413
rect -1131 1240 -1102 1413
rect -1285 1207 -1102 1240
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect -462 1270 -255 1474
rect 1139 1472 1342 1480
rect -462 1139 -407 1270
rect -294 1139 -255 1270
rect -1285 863 -1102 888
rect -1285 690 -1256 863
rect -1131 690 -1102 863
rect -1285 657 -1102 690
rect -885 863 -702 888
rect -885 690 -856 863
rect -731 690 -702 863
rect -885 657 -702 690
rect -462 679 -255 1139
rect -462 548 -407 679
rect -294 548 -255 679
rect -1285 213 -1102 238
rect -1285 40 -1256 213
rect -1131 40 -1102 213
rect -1285 7 -1102 40
rect -885 213 -702 238
rect -885 40 -856 213
rect -731 40 -702 213
rect -885 7 -702 40
rect -462 -51 -255 548
rect -462 -182 -407 -51
rect -294 -182 -255 -51
rect -462 -278 -255 -182
rect 1138 1424 1342 1472
rect 1138 1293 1193 1424
rect 1306 1293 1342 1424
rect 1138 775 1342 1293
rect 1678 1268 1857 1298
rect 1678 1148 1714 1268
rect 1826 1148 1857 1268
rect 1678 1115 1857 1148
rect 2078 1268 2257 1298
rect 2078 1148 2114 1268
rect 2226 1148 2257 1268
rect 2078 1115 2257 1148
rect 1138 644 1193 775
rect 1306 659 1342 775
rect 1305 644 1342 659
rect 1138 -55 1342 644
rect 1678 618 1857 649
rect 1678 498 1714 618
rect 1826 498 1857 618
rect 1678 465 1857 498
rect 2078 618 2257 649
rect 2078 498 2114 618
rect 2226 498 2257 618
rect 2078 465 2257 498
rect 1138 -178 1341 -55
rect 1138 -278 1342 -178
rect -462 -323 1342 -278
rect -460 -412 1342 -323
<< via3 >>
rect 1714 2607 1826 2727
rect 2114 2607 2226 2727
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect 1714 1728 1826 1848
rect 2114 1728 2226 1848
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect -1256 690 -1131 863
rect -856 690 -731 863
rect -1256 40 -1131 213
rect -856 40 -731 213
rect 1714 1148 1826 1268
rect 2114 1148 2226 1268
rect 1714 498 1826 618
rect 2114 498 2226 618
<< metal4 >>
rect 1662 2727 2269 2778
rect 1662 2675 1714 2727
rect 1664 2607 1714 2675
rect 1826 2607 2114 2727
rect 2226 2607 2269 2727
rect 1664 2527 2269 2607
rect 1663 2458 2269 2527
rect 1664 2389 2269 2458
rect -1285 2319 -1102 2342
rect -1285 2146 -1256 2319
rect -1131 2146 -1102 2319
rect -1285 2113 -1102 2146
rect -885 2319 -702 2342
rect -885 2146 -856 2319
rect -731 2146 -702 2319
rect -885 2113 -702 2146
rect 1668 1848 2266 2389
rect 1668 1728 1714 1848
rect 1826 1728 2114 1848
rect 2226 1728 2266 1848
rect -1285 1413 -1102 1438
rect -1285 1240 -1256 1413
rect -1131 1240 -1102 1413
rect -1285 1207 -1102 1240
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect 1668 1268 2266 1728
rect 1668 1148 1714 1268
rect 1826 1148 2114 1268
rect 2226 1148 2266 1268
rect -1285 863 -1102 888
rect -1285 690 -1256 863
rect -1131 690 -1102 863
rect -1285 657 -1102 690
rect -885 863 -702 888
rect -885 690 -856 863
rect -731 690 -702 863
rect -885 657 -702 690
rect 1668 618 2266 1148
rect 1668 498 1714 618
rect 1826 498 2114 618
rect 2226 498 2266 618
rect -1285 213 -1102 238
rect -1285 40 -1256 213
rect -1131 40 -1102 213
rect -1285 7 -1102 40
rect -885 213 -702 238
rect -885 40 -856 213
rect -731 40 -702 213
rect -885 7 -702 40
rect 1668 -403 2266 498
rect 1668 -437 2251 -403
<< via4 >>
rect -1256 2146 -1131 2319
rect -856 2146 -731 2319
rect -1256 1240 -1131 1413
rect -856 1240 -731 1413
rect -1256 690 -1131 863
rect -856 690 -731 863
rect -1256 40 -1131 213
rect -856 40 -731 213
<< metal5 >>
rect -1299 2536 -675 2778
rect -1296 2319 -677 2536
rect -1296 2146 -1256 2319
rect -1131 2146 -856 2319
rect -731 2146 -677 2319
rect -1296 1413 -677 2146
rect -1296 1240 -1256 1413
rect -1131 1240 -856 1413
rect -731 1240 -677 1413
rect -1296 863 -677 1240
rect -1296 690 -1256 863
rect -1131 690 -856 863
rect -731 690 -677 863
rect -1296 213 -677 690
rect -1296 40 -1256 213
rect -1131 40 -856 213
rect -731 40 -677 213
rect -1296 -442 -677 40
use SR_latch  SR_latch_0 ~/mycomparator_copy1/layout/latch
timestamp 1646810677
transform 1 0 197 0 1 2227
box 0 0 436 474
use latch_2  latch_2_0 ~/mycomparator/layout/latch
timestamp 1647337196
transform 1 0 43 0 1 1318
box 0 0 801 501
use preamp_part1  preamp_part1_0 ~/mycomparator/layout/preamp
timestamp 1646810354
transform 1 0 360 0 1 130
box -360 -130 510 508
use preamp_part2  preamp_part2_0 ~/mycomparator/layout/preamp
timestamp 1646810398
transform 1 0 69 0 1 688
box 58 1 641 544
<< labels >>
rlabel metal3 413 -412 413 -412 5 CLK
rlabel metal1 220 -58 220 -58 5 Vn
rlabel metal1 640 -58 640 -58 5 Vp
rlabel locali 257 2431 257 2431 7 Outp
rlabel locali 595 2448 595 2448 3 Outn
rlabel metal5 -988 -442 -988 -442 5 GND
rlabel metal4 2008 -437 2008 -437 5 VDD
rlabel poly 483 1945 483 1945 1 CLKBAR
<< end >>
