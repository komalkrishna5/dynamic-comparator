magic
tech sky130A
timestamp 1646832626
<< nwell >>
rect 391 2526 470 2668
rect -174 1576 74 1784
rect 89 1039 812 1201
rect 88 389 203 522
<< psubdiff >>
rect 43 64 79 76
rect 43 -12 79 0
<< nsubdiff >>
rect 405 2635 444 2647
rect 405 2533 444 2545
rect -21 1712 13 1724
rect -21 1638 13 1650
rect 166 1154 208 1166
rect 166 1069 208 1081
rect 97 504 156 516
rect 97 392 156 404
<< psubdiffcont >>
rect 43 0 79 64
<< nsubdiffcont >>
rect 405 2545 444 2635
rect -21 1650 13 1712
rect 166 1081 208 1154
rect 97 404 156 504
<< poly >>
rect 77 2461 131 2474
rect 77 2435 89 2461
rect 114 2458 131 2461
rect 114 2436 341 2458
rect 114 2435 131 2436
rect 77 2421 131 2435
rect 326 2406 341 2436
rect 684 2290 721 2300
rect 684 2289 692 2290
rect 524 2266 692 2289
rect 713 2266 721 2290
rect 684 2259 721 2266
rect 381 1528 493 1598
rect 255 1278 292 1288
rect 255 1259 265 1278
rect 283 1259 292 1278
rect 255 1247 292 1259
rect 545 1278 582 1288
rect 545 1259 555 1278
rect 573 1259 582 1278
rect 545 1247 582 1259
rect 265 1174 280 1247
rect 556 1175 571 1247
rect 409 745 424 803
rect 408 661 424 745
rect 407 638 425 661
rect 401 630 435 638
rect 401 609 409 630
rect 429 609 435 630
rect 401 600 435 609
<< polycont >>
rect 89 2435 114 2461
rect 692 2266 713 2290
rect 265 1259 283 1278
rect 555 1259 573 1278
rect 409 609 429 630
<< locali >>
rect 1738 2711 1798 2714
rect 1573 2704 1798 2711
rect 411 2643 440 2687
rect 574 2676 1798 2704
rect 1573 2671 1798 2676
rect 405 2635 444 2643
rect 405 2537 444 2545
rect 77 2461 131 2474
rect 77 2435 89 2461
rect 114 2435 131 2461
rect 77 2420 131 2435
rect 257 2426 388 2460
rect 545 2431 595 2468
rect 684 2290 721 2300
rect -558 2268 214 2275
rect -618 2208 214 2268
rect 684 2266 692 2290
rect 713 2266 721 2290
rect 684 2259 721 2266
rect 1738 2243 1798 2671
rect -885 2163 -702 2188
rect -885 1990 -856 2163
rect -731 2104 -702 2163
rect -618 2104 -542 2208
rect -731 2037 -542 2104
rect 1736 2165 1798 2243
rect -731 2029 -545 2037
rect -731 1990 -702 2029
rect -885 1957 -702 1990
rect 1736 1878 1795 2165
rect -25 1849 16 1855
rect -25 1819 -19 1849
rect 10 1819 16 1849
rect -25 1811 16 1819
rect 1678 1848 1856 1878
rect -14 1720 5 1811
rect 1678 1792 1714 1848
rect 1678 1728 1714 1767
rect 1826 1728 1856 1848
rect -21 1712 13 1720
rect 1678 1695 1856 1728
rect -21 1642 13 1650
rect 823 1514 851 1564
rect 823 1497 828 1514
rect 846 1497 851 1514
rect 823 1496 851 1497
rect -885 1413 -702 1438
rect 1159 1424 1335 1449
rect 1159 1422 1193 1424
rect -885 1240 -856 1413
rect -731 1382 -702 1413
rect 1160 1386 1193 1422
rect -731 1381 -17 1382
rect -731 1355 42 1381
rect 1159 1358 1193 1386
rect -731 1307 -701 1355
rect -16 1344 42 1355
rect -16 1318 73 1344
rect -16 1317 42 1318
rect -731 1240 -702 1307
rect -441 1270 -265 1295
rect 1160 1293 1193 1358
rect 1306 1386 1335 1424
rect 1306 1358 1337 1386
rect 1306 1293 1335 1358
rect -441 1268 -407 1270
rect -885 1207 -702 1240
rect -440 1139 -407 1268
rect -294 1139 -265 1270
rect 256 1278 291 1286
rect 256 1259 265 1278
rect 283 1259 291 1278
rect 256 1251 291 1259
rect 546 1278 581 1286
rect 546 1259 555 1278
rect 573 1259 581 1278
rect 1160 1268 1335 1293
rect 1678 1268 1856 1298
rect 546 1251 581 1259
rect 1678 1232 1714 1268
rect 40 1205 140 1232
rect 691 1231 1029 1232
rect 1641 1231 1714 1232
rect 691 1204 1714 1231
rect 1049 1203 1638 1204
rect -440 1114 -265 1139
rect 166 1154 259 1167
rect 208 1081 259 1154
rect 1678 1148 1714 1204
rect 1826 1148 1856 1268
rect 1678 1115 1856 1148
rect 166 1068 259 1081
rect -885 863 -702 888
rect -885 690 -856 863
rect -731 786 -702 863
rect -731 757 166 786
rect 1160 775 1335 800
rect -731 690 -702 757
rect -885 657 -702 690
rect -440 679 -265 704
rect -440 548 -407 679
rect -294 548 -265 679
rect 1160 666 1193 775
rect 1159 644 1193 666
rect 1306 644 1335 775
rect 401 630 435 638
rect 1159 637 1335 644
rect 401 609 409 630
rect 429 609 435 630
rect 1160 619 1335 637
rect 401 600 435 609
rect 1678 618 1856 650
rect 1678 570 1714 618
rect 825 569 1159 570
rect 1335 569 1714 570
rect -440 523 -265 548
rect -135 542 31 567
rect 825 541 1714 569
rect 97 504 213 512
rect 156 415 213 504
rect 1678 498 1714 541
rect 1826 498 1856 618
rect 1678 465 1856 498
rect 97 396 156 404
rect -885 213 -702 238
rect -885 40 -856 213
rect -731 119 -702 213
rect -731 93 13 119
rect 60 101 79 115
rect -731 40 -702 93
rect -885 7 -702 40
rect 43 64 79 101
rect 43 -8 79 0
rect -440 -51 -265 -26
rect -440 -182 -407 -51
rect -294 -75 -265 -51
rect -294 -182 -265 -161
rect -440 -208 -265 -182
<< viali >>
rect 89 2435 114 2461
rect 692 2266 713 2290
rect -856 1990 -731 2163
rect -19 1819 10 1849
rect 1714 1728 1826 1848
rect 153 1539 178 1562
rect 692 1539 717 1562
rect 828 1497 846 1514
rect -856 1240 -731 1413
rect 1193 1293 1306 1424
rect -407 1139 -294 1270
rect 265 1259 283 1278
rect 555 1259 573 1278
rect 1714 1148 1826 1268
rect -856 690 -731 863
rect -407 548 -294 679
rect 1193 644 1306 775
rect 409 609 429 630
rect 1714 498 1826 618
rect -856 40 -731 213
rect -407 -182 -294 -51
<< metal1 >>
rect 77 2469 131 2474
rect -105 2461 131 2469
rect -105 2435 89 2461
rect 114 2435 131 2461
rect -105 2427 131 2435
rect -105 2388 -63 2427
rect 77 2420 131 2427
rect -104 2340 -64 2388
rect -885 2163 -702 2188
rect -885 1990 -856 2163
rect -731 1990 -702 2163
rect -885 1957 -702 1990
rect -105 1896 -64 2340
rect 684 2290 721 2300
rect 684 2266 692 2290
rect 713 2285 986 2290
rect 713 2267 988 2285
rect 713 2266 721 2267
rect 684 2259 721 2266
rect 943 2244 988 2267
rect 945 1961 986 2244
rect -104 1564 -64 1896
rect -25 1849 16 1855
rect 402 1851 521 1864
rect 402 1849 433 1851
rect -25 1819 -19 1849
rect 10 1819 433 1849
rect -25 1818 433 1819
rect -25 1811 16 1818
rect 402 1811 433 1818
rect 485 1811 521 1851
rect 402 1800 521 1811
rect 136 1564 187 1572
rect -104 1562 187 1564
rect -104 1539 153 1562
rect 178 1539 187 1562
rect -104 1536 187 1539
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect -441 1270 -265 1295
rect -441 1139 -407 1270
rect -294 1139 -265 1270
rect -441 1114 -265 1139
rect -885 863 -702 888
rect -885 690 -856 863
rect -731 690 -702 863
rect -885 657 -702 690
rect -441 679 -265 704
rect -441 548 -407 679
rect -294 548 -265 679
rect -441 523 -265 548
rect -885 213 -702 238
rect -885 40 -856 213
rect -731 40 -702 213
rect -104 199 -64 1536
rect 136 1515 187 1536
rect 684 1562 726 1572
rect 684 1539 692 1562
rect 717 1561 726 1562
rect 946 1561 986 1961
rect 1678 1848 1857 1878
rect 1678 1728 1714 1848
rect 1826 1728 1857 1848
rect 1678 1695 1857 1728
rect 717 1539 987 1561
rect 684 1536 987 1539
rect 684 1530 726 1536
rect 823 1515 852 1520
rect 136 1514 852 1515
rect 136 1497 828 1514
rect 846 1497 852 1514
rect 946 1501 987 1536
rect 136 1496 852 1497
rect 823 1490 852 1496
rect 256 1282 291 1286
rect 256 1256 262 1282
rect 288 1256 291 1282
rect 256 1251 291 1256
rect 546 1282 581 1286
rect 546 1256 552 1282
rect 578 1256 581 1282
rect 546 1251 581 1256
rect -29 965 153 996
rect 601 969 903 1000
rect -29 293 -1 965
rect 130 950 153 965
rect 130 944 152 950
rect 401 634 435 638
rect 401 605 405 634
rect 433 605 435 634
rect 401 600 435 605
rect 875 293 903 969
rect -29 272 20 293
rect 858 272 903 293
rect 947 206 987 1501
rect 1159 1424 1335 1449
rect 1159 1293 1193 1424
rect 1306 1293 1335 1424
rect 1159 1268 1335 1293
rect 1678 1268 1857 1298
rect 1678 1148 1714 1268
rect 1826 1148 1857 1268
rect 1678 1115 1857 1148
rect 1159 775 1335 800
rect 1159 644 1193 775
rect 1306 644 1335 775
rect 1159 619 1335 644
rect 1678 618 1857 649
rect 1678 498 1714 618
rect 1826 498 1857 618
rect 1678 465 1857 498
rect -104 171 35 199
rect 819 178 987 206
rect -885 7 -702 40
rect -441 -51 -265 -26
rect -441 -182 -407 -51
rect -294 -182 -265 -51
rect 148 -58 295 54
rect 558 -58 708 56
rect -441 -208 -265 -182
<< via1 >>
rect -856 1990 -731 2163
rect 433 1811 485 1851
rect -856 1240 -731 1413
rect -407 1139 -294 1270
rect -856 690 -731 863
rect -407 548 -294 679
rect -856 40 -731 213
rect 1714 1728 1826 1848
rect 262 1278 288 1282
rect 262 1259 265 1278
rect 265 1259 283 1278
rect 283 1259 288 1278
rect 262 1256 288 1259
rect 552 1278 578 1282
rect 552 1259 555 1278
rect 555 1259 573 1278
rect 573 1259 578 1278
rect 552 1256 578 1259
rect 212 603 240 634
rect 405 630 433 634
rect 405 609 409 630
rect 409 609 429 630
rect 429 609 433 630
rect 405 605 433 609
rect 617 605 645 634
rect 1193 1293 1306 1424
rect 1714 1148 1826 1268
rect 1193 659 1306 775
rect 1193 644 1305 659
rect 1714 498 1826 618
rect -407 -182 -294 -51
rect 406 5 455 49
<< metal2 >>
rect -885 2163 -702 2188
rect -885 1990 -856 2163
rect -731 1990 -702 2163
rect -885 1957 -702 1990
rect 402 1851 516 1859
rect 402 1811 433 1851
rect 485 1843 516 1851
rect 1678 1848 1857 1878
rect 1678 1843 1714 1848
rect 485 1811 1714 1843
rect 402 1810 1714 1811
rect 402 1801 516 1810
rect 1678 1728 1714 1810
rect 1826 1728 1857 1848
rect 1678 1695 1857 1728
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect 1159 1433 1335 1449
rect 1159 1424 1337 1433
rect -885 1207 -702 1240
rect -441 1279 -265 1295
rect 1159 1293 1193 1424
rect 1306 1409 1337 1424
rect 1306 1314 1335 1409
rect 1306 1293 1334 1314
rect 1159 1290 1334 1293
rect 578 1289 1334 1290
rect 255 1282 292 1288
rect 255 1279 262 1282
rect -441 1270 262 1279
rect -441 1139 -407 1270
rect -294 1256 262 1270
rect 288 1256 292 1282
rect -294 1255 292 1256
rect -294 1139 -265 1255
rect 255 1247 292 1255
rect 545 1282 1334 1289
rect 545 1256 552 1282
rect 578 1268 1334 1282
rect 1678 1268 1857 1298
rect 578 1263 1325 1268
rect 578 1256 582 1263
rect 545 1247 582 1256
rect -441 1114 -265 1139
rect -397 1046 -308 1114
rect 1194 1048 1309 1263
rect 1678 1148 1714 1268
rect 1826 1148 1857 1268
rect 1678 1115 1857 1148
rect -397 1013 185 1046
rect 660 1016 1309 1048
rect -397 1012 -274 1013
rect 660 1012 1267 1016
rect -885 863 -702 888
rect -885 690 -856 863
rect -731 690 -702 863
rect 1159 775 1335 800
rect -885 657 -702 690
rect -441 679 -265 704
rect 1159 685 1193 775
rect -441 548 -407 679
rect -294 676 -265 679
rect 400 677 436 678
rect 206 676 436 677
rect -294 652 436 676
rect -294 548 -265 652
rect 206 634 243 652
rect 206 603 212 634
rect 240 603 243 634
rect 206 600 243 603
rect 400 634 436 652
rect 617 660 1193 685
rect 617 638 647 660
rect 400 605 405 634
rect 433 605 436 634
rect 400 600 436 605
rect 613 634 647 638
rect 613 605 617 634
rect 645 605 647 634
rect 1159 644 1193 660
rect 1306 659 1335 775
rect 1159 619 1305 644
rect 613 600 647 605
rect 1678 618 1857 649
rect -441 523 -265 548
rect 1678 498 1714 618
rect 1826 498 1857 618
rect 1678 465 1857 498
rect -885 213 -702 238
rect -885 40 -856 213
rect -731 40 -702 213
rect -885 7 -702 40
rect 397 49 464 55
rect 397 5 406 49
rect 455 5 464 49
rect -441 -51 -265 -26
rect -441 -182 -407 -51
rect -294 -105 -265 -51
rect 397 -105 464 5
rect -294 -150 465 -105
rect -294 -182 -265 -150
rect -441 -208 -265 -182
<< via2 >>
rect -856 1990 -731 2163
rect 1714 1728 1826 1848
rect -856 1240 -731 1413
rect 1193 1293 1306 1424
rect -407 1139 -294 1270
rect 1714 1148 1826 1268
rect -856 690 -731 863
rect -407 548 -294 679
rect 1193 659 1306 775
rect 1193 644 1305 659
rect 1714 498 1826 618
rect -856 40 -731 213
rect -407 -182 -294 -51
<< metal3 >>
rect -885 2163 -702 2188
rect -885 1990 -856 2163
rect -731 1990 -702 2163
rect -885 1957 -702 1990
rect 1678 1848 1857 1878
rect 1678 1728 1714 1848
rect 1826 1728 1857 1848
rect 1678 1695 1857 1728
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect -462 1270 -255 1474
rect -462 1139 -407 1270
rect -294 1139 -255 1270
rect -885 863 -702 888
rect -885 690 -856 863
rect -731 690 -702 863
rect -885 657 -702 690
rect -462 679 -255 1139
rect -462 548 -407 679
rect -294 548 -255 679
rect -885 213 -702 238
rect -885 40 -856 213
rect -731 40 -702 213
rect -885 7 -702 40
rect -462 -51 -255 548
rect -462 -182 -407 -51
rect -294 -182 -255 -51
rect -462 -278 -255 -182
rect 1138 1424 1342 1472
rect 1138 1293 1193 1424
rect 1306 1293 1342 1424
rect 1138 775 1342 1293
rect 1678 1268 1857 1298
rect 1678 1148 1714 1268
rect 1826 1148 1857 1268
rect 1678 1115 1857 1148
rect 1138 644 1193 775
rect 1306 659 1342 775
rect 1305 644 1342 659
rect 1138 -55 1342 644
rect 1678 618 1857 649
rect 1678 498 1714 618
rect 1826 498 1857 618
rect 1678 465 1857 498
rect 1138 -178 1341 -55
rect 1138 -278 1342 -178
rect -462 -323 1342 -278
rect -460 -412 1342 -323
<< via3 >>
rect -856 1990 -731 2163
rect 1714 1728 1826 1848
rect -856 1240 -731 1413
rect -856 690 -731 863
rect -856 40 -731 213
rect 1714 1148 1826 1268
rect 1714 498 1826 618
<< metal4 >>
rect -885 2163 -702 2188
rect -885 1990 -856 2163
rect -731 1990 -702 2163
rect -885 1957 -702 1990
rect 1670 1848 1864 2283
rect 1670 1728 1714 1848
rect 1826 1728 1864 1848
rect -885 1413 -702 1438
rect -885 1240 -856 1413
rect -731 1240 -702 1413
rect -885 1207 -702 1240
rect 1670 1268 1864 1728
rect 1670 1148 1714 1268
rect 1826 1148 1864 1268
rect -885 863 -702 888
rect -885 690 -856 863
rect -731 690 -702 863
rect -885 657 -702 690
rect 1670 618 1864 1148
rect 1670 498 1714 618
rect 1826 498 1864 618
rect -885 213 -702 238
rect -885 40 -856 213
rect -731 40 -702 213
rect -885 7 -702 40
rect 1670 -436 1864 498
<< via4 >>
rect -856 1990 -731 2163
rect -856 1240 -731 1413
rect -856 690 -731 863
rect -856 40 -731 213
<< metal5 >>
rect -897 2163 -666 2283
rect -897 1990 -856 2163
rect -731 1990 -666 2163
rect -897 1702 -666 1990
rect -889 1413 -679 1702
rect -889 1240 -856 1413
rect -731 1240 -679 1413
rect -889 863 -679 1240
rect -889 690 -856 863
rect -731 690 -679 863
rect -889 213 -679 690
rect -889 40 -856 213
rect -731 40 -679 213
rect -889 -436 -679 40
use SR_latch  SR_latch_0 ~/mycomparator_copy1/layout/latch
timestamp 1646810677
transform 1 0 197 0 1 2227
box 0 0 436 474
use latch_2  latch_2_0 ~/mycomparator/layout/latch
timestamp 1646831438
transform 1 0 43 0 1 1318
box 0 0 801 501
use preamp_part1  preamp_part1_0 ~/mycomparator/layout/preamp
timestamp 1646810354
transform 1 0 360 0 1 130
box -360 -130 510 508
use preamp_part2  preamp_part2_0 ~/mycomparator/layout/preamp
timestamp 1646810398
transform 1 0 69 0 1 688
box 58 1 641 544
<< labels >>
rlabel metal5 -785 -436 -785 -436 5 GND
rlabel metal3 394 -412 394 -412 5 CLK
rlabel metal4 1760 -436 1760 -436 5 VDD
rlabel metal1 215 -58 215 -58 5 Vn
rlabel metal1 633 -58 633 -58 5 Vp
rlabel poly 430 1528 430 1528 5 CLKBAR
rlabel metal1 966 2018 966 2018 1 Dn
rlabel metal1 -84 2018 -84 2018 1 Dp
rlabel locali 257 2432 257 2432 7 Outp
rlabel locali 595 2449 595 2449 3 Outn
<< end >>
