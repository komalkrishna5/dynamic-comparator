magic
tech sky130A
magscale 1 2
timestamp 1646261223
<< error_p >>
rect -737 162 833 200
rect -833 -162 833 162
rect -833 -200 737 -162
rect -637 -412 -625 -384
rect -637 -414 -607 -412
<< nwell >>
rect -737 162 833 200
rect -833 -162 833 162
rect -833 -200 737 -162
<< pmos >>
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
<< ndiff >>
rect -637 -414 -625 -412
<< pdiff >>
rect -793 74 -735 100
rect -797 62 -735 74
rect -797 -62 -785 62
rect -751 -62 -735 62
rect -797 -74 -735 -62
rect -793 -100 -735 -74
rect -705 62 -639 100
rect -705 -62 -689 62
rect -655 -62 -639 62
rect -705 -100 -639 -62
rect -609 62 -543 100
rect -609 -62 -593 62
rect -559 -62 -543 62
rect -609 -100 -543 -62
rect -513 62 -447 100
rect -513 -62 -497 62
rect -463 -62 -447 62
rect -513 -100 -447 -62
rect -417 62 -351 100
rect -417 -62 -401 62
rect -367 -62 -351 62
rect -417 -100 -351 -62
rect -321 62 -255 100
rect -321 -62 -305 62
rect -271 -62 -255 62
rect -321 -100 -255 -62
rect -225 62 -159 100
rect -225 -62 -209 62
rect -175 -62 -159 62
rect -225 -100 -159 -62
rect -129 62 -63 100
rect -129 -62 -113 62
rect -79 -62 -63 62
rect -129 -100 -63 -62
rect -33 62 33 100
rect -33 -62 -17 62
rect 17 -62 33 62
rect -33 -100 33 -62
rect 63 62 129 100
rect 63 -62 79 62
rect 113 -62 129 62
rect 63 -100 129 -62
rect 159 62 225 100
rect 159 -62 175 62
rect 209 -62 225 62
rect 159 -100 225 -62
rect 255 62 321 100
rect 255 -62 271 62
rect 305 -62 321 62
rect 255 -100 321 -62
rect 351 62 417 100
rect 351 -62 367 62
rect 401 -62 417 62
rect 351 -100 417 -62
rect 447 62 513 100
rect 447 -62 463 62
rect 497 -62 513 62
rect 447 -100 513 -62
rect 543 62 609 100
rect 543 -62 559 62
rect 593 -62 609 62
rect 543 -100 609 -62
rect 639 62 705 100
rect 639 -62 655 62
rect 689 -62 705 62
rect 639 -100 705 -62
rect 735 74 793 100
rect 735 62 797 74
rect 735 -62 751 62
rect 785 -62 797 62
rect 735 -74 797 -62
rect 735 -100 793 -74
<< pdiffc >>
rect -785 -62 -751 62
rect -689 -62 -655 62
rect -593 -62 -559 62
rect -497 -62 -463 62
rect -401 -62 -367 62
rect -305 -62 -271 62
rect -209 -62 -175 62
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
rect 175 -62 209 62
rect 271 -62 305 62
rect 367 -62 401 62
rect 463 -62 497 62
rect 559 -62 593 62
rect 655 -62 689 62
rect 751 -62 785 62
<< poly >>
rect -735 100 -705 126
rect -639 100 -609 130
rect -543 100 -513 126
rect -447 100 -417 130
rect -351 100 -321 126
rect -255 100 -225 130
rect -159 100 -129 126
rect -63 100 -33 130
rect 33 100 63 126
rect 129 100 159 130
rect 225 100 255 126
rect 321 100 351 130
rect 417 100 447 126
rect 513 100 543 130
rect 609 100 639 126
rect 705 100 735 130
rect -735 -116 -705 -100
rect -639 -116 -609 -100
rect -543 -116 -513 -100
rect -447 -116 -417 -100
rect -351 -116 -321 -100
rect -255 -116 -225 -100
rect -159 -116 -129 -100
rect -63 -116 -33 -100
rect 33 -116 63 -100
rect 129 -116 159 -100
rect 225 -116 255 -100
rect 321 -116 351 -100
rect 417 -116 447 -100
rect 513 -116 543 -100
rect 609 -116 639 -100
rect 705 -116 735 -100
rect -737 -168 735 -116
rect -603 -216 -543 -168
rect -667 -236 -543 -216
rect -667 -282 -651 -236
rect -601 -282 -543 -236
rect -667 -300 -543 -282
rect -603 -366 -543 -300
<< polycont >>
rect -651 -282 -601 -236
<< locali >>
rect -333 226 893 228
rect -883 176 893 226
rect -785 88 -751 176
rect -593 88 -559 176
rect -401 88 -367 176
rect -211 88 -177 176
rect -17 88 17 176
rect 175 88 209 176
rect 367 88 401 176
rect 559 88 593 176
rect 751 88 785 176
rect -691 -88 -689 -78
rect -211 68 -209 88
rect 497 -88 499 -84
rect 689 -88 691 -84
rect -691 -118 -655 -88
rect -497 -118 -463 -88
rect -305 -118 -271 -88
rect -113 -118 -79 -88
rect 79 -118 113 -88
rect 271 -118 305 -88
rect 463 -118 499 -88
rect 655 -118 691 -88
rect -691 -156 691 -118
rect -667 -232 -583 -216
rect -925 -236 -583 -232
rect -925 -282 -651 -236
rect -601 -282 -583 -236
rect -925 -288 -583 -282
rect -667 -300 -583 -288
rect -63 -232 25 -156
rect -63 -288 869 -232
rect -63 -340 25 -288
rect -637 -374 25 -340
rect -637 -376 -23 -374
rect -637 -414 -603 -376
rect -445 -424 -409 -376
rect -255 -422 -219 -376
rect -61 -416 -25 -376
rect -733 -698 -699 -556
rect -541 -684 -507 -542
rect -349 -688 -315 -546
rect -155 -694 -121 -552
rect 35 -698 69 -556
<< viali >>
rect -785 62 -751 88
rect -785 -62 -751 62
rect -785 -88 -751 -62
rect -689 62 -655 88
rect -689 -62 -655 62
rect -689 -88 -655 -62
rect -593 62 -559 88
rect -593 -62 -559 62
rect -593 -88 -559 -62
rect -497 62 -463 88
rect -497 -62 -463 62
rect -497 -88 -463 -62
rect -401 62 -367 88
rect -401 -62 -367 62
rect -401 -88 -367 -62
rect -305 62 -271 88
rect -305 -62 -271 62
rect -305 -88 -271 -62
rect -209 62 -175 88
rect -209 -62 -175 62
rect -209 -88 -175 -62
rect -113 62 -79 88
rect -113 -62 -79 62
rect -113 -88 -79 -62
rect -17 62 17 88
rect -17 -62 17 62
rect -17 -88 17 -62
rect 79 62 113 88
rect 79 -62 113 62
rect 79 -88 113 -62
rect 175 62 209 88
rect 175 -62 209 62
rect 175 -88 209 -62
rect 271 62 305 88
rect 271 -62 305 62
rect 271 -88 305 -62
rect 367 62 401 88
rect 367 -62 401 62
rect 367 -88 401 -62
rect 463 62 497 88
rect 463 -62 497 62
rect 463 -88 497 -62
rect 559 62 593 88
rect 559 -62 593 62
rect 559 -88 593 -62
rect 655 62 689 88
rect 655 -62 689 62
rect 655 -88 689 -62
rect 751 62 785 88
rect 751 -62 785 62
rect 751 -88 785 -62
<< metal1 >>
rect -791 88 -745 100
rect -791 -88 -785 88
rect -751 -88 -745 88
rect -791 -100 -745 -88
rect -695 88 -649 100
rect -695 -88 -689 88
rect -655 -88 -649 88
rect -695 -100 -649 -88
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -503 88 -457 100
rect -503 -88 -497 88
rect -463 -88 -457 88
rect -503 -100 -457 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 457 88 503 100
rect 457 -88 463 88
rect 497 -88 503 88
rect 457 -100 503 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
rect 649 88 695 100
rect 649 -88 655 88
rect 689 -88 695 88
rect 649 -100 695 -88
rect 745 88 791 100
rect 745 -88 751 88
rect 785 -88 791 88
rect 745 -100 791 -88
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 16 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
