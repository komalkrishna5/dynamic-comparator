magic
tech sky130A
magscale 1 2
timestamp 1646810591
<< locali >>
rect 502 900 1140 950
rect 628 796 662 900
rect 820 802 854 900
rect 480 436 1120 492
rect 520 0 1092 52
<< metal1 >>
rect 718 962 956 1002
rect 718 782 764 962
rect 910 784 956 962
use inv_W2  inv_W2_0 ~/mycomparator/layout/myinv_layout2
timestamp 1646730554
transform 1 0 120 0 1 72
box -120 -72 404 878
use inv_W2  inv_W2_1
timestamp 1646730554
transform 1 0 1198 0 1 72
box -120 -72 404 878
use sky130_fd_pr__pfet_01v8_5SVZDE  sky130_fd_pr__pfet_01v8_5SVZDE_0
timestamp 1646503715
transform 1 0 789 0 1 712
box -789 -196 805 222
<< labels >>
rlabel space 1602 26 1602 26 3 GND
rlabel space 1602 936 1602 936 3 VDD
<< end >>
