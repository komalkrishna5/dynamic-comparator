magic
tech sky130A
timestamp 1645264122
<< locali >>
rect -1 451 17 475
rect 0 218 21 246
rect 475 218 488 246
rect 0 1 22 27
use inv_W1  inv_W1_0
timestamp 1645263751
transform 1 0 50 0 1 36
box -50 -36 194 439
use inv_W1  inv_W1_1
timestamp 1645263751
transform 1 0 294 0 1 36
box -50 -36 194 439
<< labels >>
rlabel locali 0 6 0 6 7 GND
rlabel locali 0 227 0 227 7 Vin
rlabel locali -1 456 -1 456 7 VDD
rlabel locali 488 227 488 227 3 Vout
<< end >>
