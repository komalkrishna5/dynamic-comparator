* SPICE3 file created from comparator_v3.ext - technology: sky130A

.subckt sky130_fd_pr__diode_pw2nd_05v5_KLAK3C a_n45_n45# w_n183_n183#
D0 w_n183_n183# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
.ends

.subckt sky130_fd_pr__pfet_01v8_RFM3CD a_n73_n100# w_n109_n162# a_15_n100# a_n15_n126#
+ VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# w_n109_n162# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_F5U58G#0 a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_XJTKXQ#0 a_n63_n152# a_63_n100# a_n125_n74# a_n33_n100#
+ VSUBS
X0 a_63_n100# a_n63_n152# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n152# a_n125_n74# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt preamp_part2 a_148_644# sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126# a_380_480#
+ sky130_fd_pr__pfet_01v8_RFM3CD_1/w_n109_n162# sky130_fd_pr__pfet_01v8_RFM3CD_0/a_n15_n126#
+ sky130_fd_pr__pfet_01v8_RFM3CD_1/a_n15_n126# a_1170_652# sky130_fd_pr__pfet_01v8_RFM3CD_0/w_n109_n162#
+ VDD GND a_792_2# VSUBS
Xsky130_fd_pr__pfet_01v8_RFM3CD_0 VDD sky130_fd_pr__pfet_01v8_RFM3CD_0/w_n109_n162#
+ li_210_488# sky130_fd_pr__pfet_01v8_RFM3CD_0/a_n15_n126# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD
Xsky130_fd_pr__pfet_01v8_RFM3CD_1 li_928_394# sky130_fd_pr__pfet_01v8_RFM3CD_1/w_n109_n162#
+ VDD sky130_fd_pr__pfet_01v8_RFM3CD_1/a_n15_n126# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD
Xsky130_fd_pr__nfet_01v8_F5U58G_0 m1_322_206# GND sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126#
+ VSUBS sky130_fd_pr__nfet_01v8_F5U58G#0
Xsky130_fd_pr__nfet_01v8_F5U58G_1 a_792_2# li_210_488# a_148_644# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#0
Xsky130_fd_pr__nfet_01v8_F5U58G_2 li_928_394# a_380_480# a_1170_652# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#0
Xsky130_fd_pr__nfet_01v8_XJTKXQ_0 a_380_480# m1_322_206# m1_322_206# li_210_488# VSUBS
+ sky130_fd_pr__nfet_01v8_XJTKXQ#0
Xsky130_fd_pr__nfet_01v8_XJTKXQ_1 a_792_2# m1_322_206# m1_322_206# li_928_394# VSUBS
+ sky130_fd_pr__nfet_01v8_XJTKXQ#0
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT7GK8 a_n45_n45# w_n183_n183#
D0 w_n183_n183# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
.ends

.subckt sky130_fd_pr__nfet_01v8_F5U58G a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_AC5E9B w_n161_n200# a_33_n126# a_63_n100# a_n125_n74#
+ a_n33_n100# a_n63_n130# VSUBS
X0 a_63_n100# a_33_n126# a_n33_n100# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n130# a_n125_n74# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt SR_latch a_648_848# sky130_fd_pr__nfet_01v8_F5U58G_1/a_n15_n126# sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126#
+ a_262_508# VDD w_0_524# GND VSUBS
Xsky130_fd_pr__nfet_01v8_F5U58G_0 a_648_848# GND sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126#
+ VSUBS sky130_fd_pr__nfet_01v8_F5U58G
Xsky130_fd_pr__nfet_01v8_F5U58G_1 GND a_262_508# sky130_fd_pr__nfet_01v8_F5U58G_1/a_n15_n126#
+ VSUBS sky130_fd_pr__nfet_01v8_F5U58G
Xsky130_fd_pr__pfet_01v8_AC5E9B_0 w_0_524# a_262_508# VDD VDD a_648_848# a_262_508#
+ VSUBS sky130_fd_pr__pfet_01v8_AC5E9B
Xsky130_fd_pr__pfet_01v8_AC5E9B_1 w_0_524# a_648_848# VDD VDD a_262_508# a_648_848#
+ VSUBS sky130_fd_pr__pfet_01v8_AC5E9B
.ends

.subckt sky130_fd_pr__nfet_01v8_G6PLX8 a_159_n100# a_n221_n74# a_n129_n100# a_63_n100#
+ a_n33_n100# a_n159_n122# VSUBS
X0 a_n129_n100# a_n159_n122# a_n221_n74# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
X1 a_63_n100# a_n159_n122# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_n33_n100# a_n159_n122# a_n129_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_159_n100# a_n159_n122# a_63_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_F5U58G#1 a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_8FHE5N a_n33_n50# a_63_n50# a_n63_n76# a_33_n76# a_n125_n39#
+ VSUBS
X0 a_n33_n50# a_n63_n76# a_n125_n39# VSUBS sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.66e+06u as=1.528e+11p ps=1.62e+06u w=500000u l=150000u
X1 a_63_n50# a_33_n76# a_n33_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=1.528e+11p pd=1.62e+06u as=0p ps=0u w=500000u l=150000u
.ends

.subckt preamp_part1 li_954_42# li_n718_44# a_n656_268# a_80_n258# a_n302_940# w_n720_482#
+ a_n434_n260# a_506_940# a_864_270# VDD a_388_n260# GND VSUBS
Xsky130_fd_pr__nfet_01v8_G6PLX8_0 li_n484_188# li_n484_188# a_n656_268# a_n656_268#
+ li_n484_188# a_n434_n260# VSUBS sky130_fd_pr__nfet_01v8_G6PLX8
Xsky130_fd_pr__nfet_01v8_G6PLX8_1 li_n484_188# li_n484_188# a_864_270# a_864_270#
+ li_n484_188# a_388_n260# VSUBS sky130_fd_pr__nfet_01v8_G6PLX8
Xsky130_fd_pr__pfet_01v8_RFM3CD_0 VDD w_n720_482# a_n656_268# a_n302_940# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD
Xsky130_fd_pr__pfet_01v8_RFM3CD_1 a_864_270# w_n720_482# VDD a_506_940# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD
Xsky130_fd_pr__nfet_01v8_F5U58G_0 li_n718_44# GND a_n656_268# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#1
Xsky130_fd_pr__nfet_01v8_F5U58G_1 GND li_954_42# a_864_270# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#1
Xsky130_fd_pr__nfet_01v8_8FHE5N_0 li_n484_188# GND a_80_n258# a_80_n258# GND VSUBS
+ sky130_fd_pr__nfet_01v8_8FHE5N
.ends

.subckt sky130_fd_pr__nfet_01v8_7RYEVP a_n73_n69# a_n33_n157# a_15_n69# VSUBS
X0 a_15_n69# a_n33_n157# a_n73_n69# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt nmos_1u sky130_fd_pr__nfet_01v8_7RYEVP_0/VSUBS sky130_fd_pr__nfet_01v8_7RYEVP_0/a_15_n69#
+ m1_n86_2#
Xsky130_fd_pr__nfet_01v8_7RYEVP_0 sky130_fd_pr__nfet_01v8_7RYEVP_0/VSUBS m1_n86_2#
+ sky130_fd_pr__nfet_01v8_7RYEVP_0/a_15_n69# sky130_fd_pr__nfet_01v8_7RYEVP_0/VSUBS
+ sky130_fd_pr__nfet_01v8_7RYEVP
.ends

.subckt pmos_2uf2 a_63_n100# a_33_n130# w_n317_n202# a_n33_n100# a_n63_n130# VSUBS
X0 a_63_n100# a_33_n130# a_n33_n100# w_n317_n202# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n130# w_n317_n202# w_n317_n202# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.8e+11p ps=2.76e+06u w=1e+06u l=150000u
.ends

.subckt inv_W1 Vout Vin VDD GND
Xnmos_1u_0 GND Vout Vin nmos_1u
Xpmos_2uf2_0 VDD Vin VDD Vout Vin GND pmos_2uf2
.ends

.subckt sky130_fd_pr__pfet_01v8_AC5Z8B a_159_n100# li_217_n290# li_n261_n290# li_229_174#
+ a_n221_n74# a_n129_n100# a_n159_n152# li_225_n726# a_n33_n100# w_n261_n210# li_n261_174#
+ li_n261_n726# VSUBS
X0 a_n129_n100# a_n159_n152# a_n33_n100# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=5.32e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n159_n152# a_n129_n100# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_159_n100# a_n159_n152# a_n129_n100# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_n129_n100# a_n159_n152# a_n221_n74# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_XJTKXQ a_33_n122# a_n63_n122# a_63_n100# a_n125_n74#
+ a_n33_n100# VSUBS
X0 a_63_n100# a_33_n122# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n122# a_n125_n74# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt inv_W2 sky130_fd_pr__pfet_01v8_AC5Z8B_0/w_n261_n210# li_202_260# li_n100_828#
+ li_n100_n72# a_84_352# VSUBS
Xsky130_fd_pr__pfet_01v8_AC5Z8B_0 li_n100_828# li_202_260# a_84_352# li_n100_828#
+ li_n100_828# li_202_260# a_84_352# li_n100_n72# li_n100_828# sky130_fd_pr__pfet_01v8_AC5Z8B_0/w_n261_n210#
+ li_n100_828# li_n100_n72# VSUBS sky130_fd_pr__pfet_01v8_AC5Z8B
Xsky130_fd_pr__nfet_01v8_XJTKXQ_0 a_84_352# a_84_352# li_n100_n72# li_n100_n72# li_202_260#
+ VSUBS sky130_fd_pr__nfet_01v8_XJTKXQ
.ends

.subckt sky130_fd_pr__pfet_01v8_5SVZDE a_n111_n158# a_n173_n100# a_15_n100# a_111_n100#
+ a_n81_n100# w_n789_n196# VSUBS
X0 a_15_n100# a_n111_n158# a_n81_n100# w_n789_n196# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_111_n100# a_n111_n158# a_15_n100# w_n789_n196# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_n81_n100# a_n111_n158# a_n173_n100# w_n789_n196# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt latch_2 m1_718_782# inv_W2_1/li_202_260# li_480_436# sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196#
+ li_520_0# sky130_fd_pr__pfet_01v8_5SVZDE_0/a_n111_n158# VSUBS inv_W2_0/a_84_352#
Xinv_W2_0 sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196# li_480_436# li_502_900# li_520_0#
+ inv_W2_0/a_84_352# VSUBS inv_W2
Xinv_W2_1 sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196# inv_W2_1/li_202_260# li_502_900#
+ li_520_0# li_480_436# VSUBS inv_W2
Xsky130_fd_pr__pfet_01v8_5SVZDE_0 sky130_fd_pr__pfet_01v8_5SVZDE_0/a_n111_n158# li_502_900#
+ li_502_900# m1_718_782# m1_718_782# sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196#
+ VSUBS sky130_fd_pr__pfet_01v8_5SVZDE
C0 sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196# VSUBS 2.01fF
.ends


* Top level circuit comparator_v3

Xsky130_fd_pr__diode_pw2nd_05v5_KLAK3C_2 VDD VDD sky130_fd_pr__diode_pw2nd_05v5_KLAK3C
Xsky130_fd_pr__diode_pw2nd_05v5_KLAK3C_3 VDD VDD sky130_fd_pr__diode_pw2nd_05v5_KLAK3C
Xpreamp_part2_0 CLK CLK m1_1202_1938# VDD CLK CLK CLK VDD VDD VDD m1_n58_544# VDD
+ preamp_part2
Xsky130_fd_pr__diode_pw2nd_05v5_FT7GK8_0 VDD VDD sky130_fd_pr__diode_pw2nd_05v5_FT7GK8
Xsky130_fd_pr__diode_pw2nd_05v5_FT7GK8_1 VDD VDD sky130_fd_pr__diode_pw2nd_05v5_FT7GK8
Xsky130_fd_pr__diode_pw2nd_05v5_FT7GK8_2 VDD VDD sky130_fd_pr__diode_pw2nd_05v5_FT7GK8
Xsky130_fd_pr__diode_pw2nd_05v5_FT7GK8_3 VDD VDD sky130_fd_pr__diode_pw2nd_05v5_FT7GK8
XSR_latch_0 Outp a_1048_4532# a_154_4842# Outn VDD VDD VDD VDD SR_latch
Xpreamp_part1_0 a_1048_4532# a_154_4842# m1_n58_544# CLK CLK VDD Vn CLK m1_1202_1938#
+ VDD Vp VDD VDD preamp_part1
Xinv_W1_0 inv_W1_0/Vout CLK VDD VDD inv_W1
Xlatch_2_0 VDD a_154_4842# a_1048_4532# VDD VDD inv_W1_0/Vout VDD a_154_4842# latch_2
Xsky130_fd_pr__diode_pw2nd_05v5_KLAK3C_0 VDD VDD sky130_fd_pr__diode_pw2nd_05v5_KLAK3C
Xsky130_fd_pr__diode_pw2nd_05v5_KLAK3C_1 VDD VDD sky130_fd_pr__diode_pw2nd_05v5_KLAK3C
C0 a_1048_4532# VDD 3.13fF
C1 a_154_4842# VDD 4.97fF
C2 inv_W1_0/Vout VDD 2.30fF
C3 CLK VDD 20.76fF
C4 m1_n58_544# VDD 2.18fF
.end

