magic
tech sky130A
magscale 1 2
timestamp 1646248588
<< error_p >>
rect 19 272 77 278
rect 19 238 31 272
rect 19 232 77 238
rect -77 -238 -19 -232
rect -77 -272 -65 -238
rect -77 -278 -19 -272
<< pwell >>
rect -263 -410 263 410
<< nmos >>
rect -63 -200 -33 200
rect 33 -200 63 200
<< ndiff >>
rect -121 144 -63 200
rect -125 132 -63 144
rect -125 -132 -113 132
rect -79 -132 -63 132
rect -125 -144 -63 -132
rect -121 -200 -63 -144
rect -33 132 33 200
rect -33 -132 -17 132
rect 17 -132 33 132
rect -33 -200 33 -132
rect 63 144 121 200
rect 63 132 125 144
rect 63 -132 79 132
rect 113 -132 125 132
rect 63 -144 125 -132
rect 63 -200 121 -144
<< ndiffc >>
rect -113 -132 -79 132
rect -17 -132 17 132
rect 79 -132 113 132
<< psubdiff >>
rect -227 340 -92 374
rect 92 340 227 374
rect -227 195 -193 340
rect -227 -340 -193 -195
rect 193 195 227 340
rect 193 -340 227 -195
rect -227 -374 -92 -340
rect 92 -374 227 -340
<< psubdiffcont >>
rect -92 340 92 374
rect -227 -195 -193 195
rect 193 -195 227 195
rect -92 -374 92 -340
<< poly >>
rect 15 272 81 288
rect 15 238 31 272
rect 65 238 81 272
rect -63 200 -33 226
rect 15 222 81 238
rect 33 200 63 222
rect -63 -222 -33 -200
rect -81 -238 -15 -222
rect 33 -226 63 -200
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect -81 -288 -15 -272
<< polycont >>
rect 31 238 65 272
rect -65 -272 -31 -238
<< locali >>
rect -227 340 -92 374
rect 92 340 227 374
rect -227 195 -193 340
rect 15 238 31 272
rect 65 238 81 272
rect 193 195 227 340
rect -113 132 -79 148
rect -113 -148 -79 -132
rect -17 132 17 148
rect -17 -148 17 -132
rect 79 132 113 148
rect 79 -148 113 -132
rect -227 -340 -193 -195
rect -81 -272 -65 -238
rect -31 -272 -15 -238
rect 193 -340 227 -195
rect -227 -374 -92 -340
rect 92 -374 227 -340
<< viali >>
rect 31 238 65 272
rect -113 -132 -79 132
rect -17 -132 17 132
rect 79 -132 113 132
rect -65 -272 -31 -238
<< metal1 >>
rect 19 272 77 278
rect 19 238 31 272
rect 65 238 77 272
rect 19 232 77 238
rect -119 132 -73 144
rect -119 -132 -113 132
rect -79 -132 -73 132
rect -119 -144 -73 -132
rect -23 132 23 144
rect -23 -132 -17 132
rect 17 -132 23 132
rect -23 -144 23 -132
rect 73 132 119 144
rect 73 -132 79 132
rect 113 -132 119 132
rect 73 -144 119 -132
rect -77 -238 -19 -232
rect -77 -272 -65 -238
rect -31 -272 -19 -238
rect -77 -278 -19 -272
<< properties >>
string FIXED_BBOX -210 -357 210 357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.150 m 1 nf 2 diffcov 70 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
