magic
tech sky130A
magscale 1 2
timestamp 1646431323
<< nmos >>
rect -15 -100 15 100
<< ndiff >>
rect -73 62 -15 100
rect -73 -62 -61 62
rect -27 -62 -15 62
rect -73 -100 -15 -62
rect 15 62 73 100
rect 15 -62 27 62
rect 61 -62 73 62
rect 15 -100 73 -62
<< ndiffc >>
rect -61 -62 -27 62
rect 27 -62 61 62
<< poly >>
rect -15 100 15 126
rect -15 -126 15 -100
<< locali >>
rect -61 62 -27 78
rect -61 -78 -27 -62
rect 27 62 61 78
rect 27 -78 61 -62
<< viali >>
rect -61 -62 -27 62
rect 27 -62 61 62
<< metal1 >>
rect -67 62 -21 74
rect -67 -62 -61 62
rect -27 -62 -21 62
rect -67 -74 -21 -62
rect 21 62 67 74
rect 21 -62 27 62
rect 61 -62 67 62
rect 21 -74 67 -62
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 1 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
