magic
tech sky130A
magscale 1 2
timestamp 1646734260
<< poly >>
rect 148 706 230 722
rect 148 660 164 706
rect 214 660 230 706
rect 148 644 230 660
rect 1170 704 1246 714
rect 1170 668 1188 704
rect 1228 668 1246 704
rect 1170 652 1246 668
rect 174 576 204 644
rect 380 608 614 620
rect 380 546 536 608
rect 598 546 614 608
rect 1194 580 1224 652
rect 380 530 614 546
rect 380 480 506 530
rect 890 92 1016 226
rect 792 80 1016 92
rect 792 18 808 80
rect 870 18 1016 80
rect 792 2 1016 18
<< polycont >>
rect 164 660 214 706
rect 1188 668 1228 704
rect 536 546 598 608
rect 808 18 870 80
<< locali >>
rect 116 1034 1282 1088
rect 346 938 380 1034
rect 1016 932 1050 1034
rect 148 706 230 722
rect 148 660 164 706
rect 214 660 230 706
rect 148 644 230 660
rect 434 538 468 796
rect 210 488 468 538
rect 520 608 614 624
rect 520 546 536 608
rect 598 546 614 608
rect 520 530 614 546
rect 928 532 962 790
rect 1170 704 1246 714
rect 1170 668 1188 704
rect 1228 668 1246 704
rect 1170 652 1246 668
rect 420 396 468 488
rect 928 484 1188 532
rect 928 394 976 484
rect 722 196 756 270
rect 116 138 1282 196
rect 792 80 886 96
rect 792 18 808 80
rect 870 18 886 80
rect 792 2 886 18
<< viali >>
rect 164 660 214 706
rect 536 546 598 608
rect 1188 668 1228 704
rect 808 18 870 80
<< metal1 >>
rect 148 712 230 722
rect 148 654 158 712
rect 220 654 230 712
rect 148 644 230 654
rect 1170 710 1246 714
rect 1170 658 1180 710
rect 1236 658 1246 710
rect 1170 652 1246 658
rect 520 608 1276 624
rect 520 546 536 608
rect 598 562 1276 608
rect 598 546 614 562
rect 520 530 614 546
rect 1230 520 1276 562
rect 122 92 168 398
rect 322 244 370 288
rect 516 244 562 284
rect 628 244 674 292
rect 834 244 880 296
rect 1026 244 1072 284
rect 322 206 1072 244
rect 792 92 886 96
rect 122 80 886 92
rect 122 30 808 80
rect 792 18 808 30
rect 870 18 886 80
rect 792 2 886 18
<< via1 >>
rect 158 706 220 712
rect 158 660 164 706
rect 164 660 214 706
rect 214 660 220 706
rect 158 654 220 660
rect 1180 704 1236 710
rect 1180 668 1188 704
rect 1188 668 1228 704
rect 1228 668 1236 704
rect 1180 658 1236 668
<< metal2 >>
rect 148 714 230 722
rect 1180 714 1236 720
rect 148 712 1246 714
rect 148 654 158 712
rect 220 710 1246 712
rect 220 658 1180 710
rect 1236 658 1246 710
rect 220 654 1246 658
rect 148 652 1246 654
rect 148 644 230 652
rect 1180 648 1236 652
use sky130_fd_pr__nfet_01v8_F5U58G#0#0  sky130_fd_pr__nfet_01v8_F5U58G_0
timestamp 1646431323
transform 1 0 695 0 1 346
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_F5U58G#0#0  sky130_fd_pr__nfet_01v8_F5U58G_1
timestamp 1646431323
transform 1 0 189 0 1 458
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_F5U58G#0#0  sky130_fd_pr__nfet_01v8_F5U58G_2
timestamp 1646431323
transform 1 0 1209 0 1 460
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_XJTKXQ#0#0  sky130_fd_pr__nfet_01v8_XJTKXQ_0
timestamp 1646429429
transform 1 0 443 0 1 346
box -125 -152 125 154
use sky130_fd_pr__nfet_01v8_XJTKXQ#0#0  sky130_fd_pr__nfet_01v8_XJTKXQ_1
timestamp 1646429429
transform 1 0 953 0 1 346
box -125 -152 125 154
use sky130_fd_pr__pfet_01v8_RFM3CD#0  sky130_fd_pr__pfet_01v8_RFM3CD_0
timestamp 1646431323
transform 1 0 407 0 1 864
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_RFM3CD#0  sky130_fd_pr__pfet_01v8_RFM3CD_1
timestamp 1646431323
transform 1 0 989 0 1 864
box -109 -162 109 162
<< end >>
