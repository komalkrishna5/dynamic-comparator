magic
tech sky130A
magscale 1 2
timestamp 1646319668
<< nwell >>
rect -737 162 833 200
rect -833 -162 833 162
rect -833 -200 737 -162
<< pmos >>
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
<< pdiff >>
rect -793 74 -735 100
rect -797 62 -735 74
rect -797 -62 -785 62
rect -751 -62 -735 62
rect -797 -74 -735 -62
rect -793 -100 -735 -74
rect -705 62 -639 100
rect -705 -62 -689 62
rect -655 -62 -639 62
rect -705 -100 -639 -62
rect -609 62 -543 100
rect -609 -62 -593 62
rect -559 -62 -543 62
rect -609 -100 -543 -62
rect -513 62 -447 100
rect -513 -62 -497 62
rect -463 -62 -447 62
rect -513 -100 -447 -62
rect -417 62 -351 100
rect -417 -62 -401 62
rect -367 -62 -351 62
rect -417 -100 -351 -62
rect -321 62 -255 100
rect -321 -62 -305 62
rect -271 -62 -255 62
rect -321 -100 -255 -62
rect -225 62 -159 100
rect -225 -62 -209 62
rect -175 -62 -159 62
rect -225 -100 -159 -62
rect -129 62 -63 100
rect -129 -62 -113 62
rect -79 -62 -63 62
rect -129 -100 -63 -62
rect -33 62 33 100
rect -33 -62 -17 62
rect 17 -62 33 62
rect -33 -100 33 -62
rect 63 62 129 100
rect 63 -62 79 62
rect 113 -62 129 62
rect 63 -100 129 -62
rect 159 62 225 100
rect 159 -62 175 62
rect 209 -62 225 62
rect 159 -100 225 -62
rect 255 62 321 100
rect 255 -62 271 62
rect 305 -62 321 62
rect 255 -100 321 -62
rect 351 62 417 100
rect 351 -62 367 62
rect 401 -62 417 62
rect 351 -100 417 -62
rect 447 62 513 100
rect 447 -62 463 62
rect 497 -62 513 62
rect 447 -100 513 -62
rect 543 62 609 100
rect 543 -62 559 62
rect 593 -62 609 62
rect 543 -100 609 -62
rect 639 62 705 100
rect 639 -62 655 62
rect 689 -62 705 62
rect 639 -100 705 -62
rect 735 74 793 100
rect 735 62 797 74
rect 735 -62 751 62
rect 785 -62 797 62
rect 735 -74 797 -62
rect 735 -100 793 -74
<< pdiffc >>
rect -785 -62 -751 62
rect -689 -62 -655 62
rect -593 -62 -559 62
rect -497 -62 -463 62
rect -401 -62 -367 62
rect -305 -62 -271 62
rect -209 -62 -175 62
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
rect 175 -62 209 62
rect 271 -62 305 62
rect 367 -62 401 62
rect 463 -62 497 62
rect 559 -62 593 62
rect 655 -62 689 62
rect 751 -62 785 62
<< poly >>
rect -735 100 -705 126
rect -639 100 -609 130
rect -543 100 -513 126
rect -447 100 -417 130
rect -351 100 -321 126
rect -255 100 -225 130
rect -159 100 -129 126
rect -63 100 -33 130
rect 33 100 63 126
rect 129 100 159 130
rect 225 100 255 126
rect 321 100 351 130
rect 417 100 447 126
rect 513 100 543 130
rect 609 100 639 126
rect 705 100 735 130
rect -735 -128 -705 -100
rect -639 -126 -609 -100
rect -543 -128 -513 -100
rect -447 -126 -417 -100
rect -351 -128 -321 -100
rect -255 -126 -225 -100
rect -159 -128 -129 -100
rect -63 -126 -33 -100
rect 33 -128 63 -100
rect 129 -126 159 -100
rect 225 -128 255 -100
rect 321 -126 351 -100
rect 417 -128 447 -100
rect 513 -126 543 -100
rect 609 -128 639 -100
rect 705 -126 735 -100
<< locali >>
rect -785 62 -751 78
rect -785 -78 -751 -62
rect -689 62 -655 78
rect -689 -78 -655 -62
rect -593 62 -559 78
rect -593 -78 -559 -62
rect -497 62 -463 78
rect -497 -78 -463 -62
rect -401 62 -367 78
rect -401 -78 -367 -62
rect -305 62 -271 78
rect -305 -78 -271 -62
rect -209 62 -175 78
rect -209 -78 -175 -62
rect -113 62 -79 78
rect -113 -78 -79 -62
rect -17 62 17 78
rect -17 -78 17 -62
rect 79 62 113 78
rect 79 -78 113 -62
rect 175 62 209 78
rect 175 -78 209 -62
rect 271 62 305 78
rect 271 -78 305 -62
rect 367 62 401 78
rect 367 -78 401 -62
rect 463 62 497 78
rect 463 -78 497 -62
rect 559 62 593 78
rect 559 -78 593 -62
rect 655 62 689 78
rect 655 -78 689 -62
rect 751 62 785 78
rect 751 -78 785 -62
<< viali >>
rect -785 -62 -751 62
rect -689 -62 -655 62
rect -593 -62 -559 62
rect -497 -62 -463 62
rect -401 -62 -367 62
rect -305 -62 -271 62
rect -209 -62 -175 62
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
rect 175 -62 209 62
rect 271 -62 305 62
rect 367 -62 401 62
rect 463 -62 497 62
rect 559 -62 593 62
rect 655 -62 689 62
rect 751 -62 785 62
<< metal1 >>
rect -791 62 -745 74
rect -791 -62 -785 62
rect -751 -62 -745 62
rect -791 -74 -745 -62
rect -695 62 -649 74
rect -695 -62 -689 62
rect -655 -62 -649 62
rect -695 -74 -649 -62
rect -599 62 -553 74
rect -599 -62 -593 62
rect -559 -62 -553 62
rect -599 -74 -553 -62
rect -503 62 -457 74
rect -503 -62 -497 62
rect -463 -62 -457 62
rect -503 -74 -457 -62
rect -407 62 -361 74
rect -407 -62 -401 62
rect -367 -62 -361 62
rect -407 -74 -361 -62
rect -311 62 -265 74
rect -311 -62 -305 62
rect -271 -62 -265 62
rect -311 -74 -265 -62
rect -215 62 -169 74
rect -215 -62 -209 62
rect -175 -62 -169 62
rect -215 -74 -169 -62
rect -119 62 -73 74
rect -119 -62 -113 62
rect -79 -62 -73 62
rect -119 -74 -73 -62
rect -23 62 23 74
rect -23 -62 -17 62
rect 17 -62 23 62
rect -23 -74 23 -62
rect 73 62 119 74
rect 73 -62 79 62
rect 113 -62 119 62
rect 73 -74 119 -62
rect 169 62 215 74
rect 169 -62 175 62
rect 209 -62 215 62
rect 169 -74 215 -62
rect 265 62 311 74
rect 265 -62 271 62
rect 305 -62 311 62
rect 265 -74 311 -62
rect 361 62 407 74
rect 361 -62 367 62
rect 401 -62 407 62
rect 361 -74 407 -62
rect 457 62 503 74
rect 457 -62 463 62
rect 497 -62 503 62
rect 457 -74 503 -62
rect 553 62 599 74
rect 553 -62 559 62
rect 593 -62 599 62
rect 553 -74 599 -62
rect 649 62 695 74
rect 649 -62 655 62
rect 689 -62 695 62
rect 649 -74 695 -62
rect 745 62 791 74
rect 745 -62 751 62
rect 785 -62 791 62
rect 745 -74 791 -62
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 16 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
