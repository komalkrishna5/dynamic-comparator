magic
tech sky130A
magscale 1 2
timestamp 1646734260
<< nwell >>
rect -720 482 1018 816
<< poly >>
rect -302 1000 -234 1016
rect -302 958 -286 1000
rect -250 958 -234 1000
rect -302 940 -234 958
rect 506 1000 574 1016
rect 506 958 522 1000
rect 562 958 574 1000
rect 506 940 574 958
rect -282 754 -252 940
rect 524 764 556 940
rect -656 326 -594 342
rect -656 284 -640 326
rect -606 284 -594 326
rect -656 268 -594 284
rect 864 328 926 344
rect 864 286 880 328
rect 914 286 926 328
rect 864 270 926 286
rect -640 242 -610 268
rect 882 234 912 270
rect -434 4 -404 6
rect -338 4 -308 6
rect -242 4 -212 6
rect -146 4 -116 6
rect -434 -168 -116 4
rect -434 -234 -406 -168
rect -144 -234 -116 -168
rect -434 -260 -116 -234
rect 80 -170 206 58
rect 80 -238 104 -170
rect 180 -238 206 -170
rect 80 -258 206 -238
rect 388 -2 418 4
rect 484 -2 514 4
rect 580 -2 610 4
rect 676 -2 706 4
rect 388 -164 706 -2
rect 388 -234 414 -164
rect 680 -234 706 -164
rect 388 -260 706 -234
<< polycont >>
rect -286 958 -250 1000
rect 522 958 562 1000
rect -640 284 -606 326
rect 880 286 914 328
rect -406 -234 -144 -168
rect 104 -238 180 -170
rect 414 -234 680 -164
<< locali >>
rect -302 1000 -234 1016
rect -302 958 -286 1000
rect -250 958 -234 1000
rect -302 940 -234 958
rect 506 1000 574 1016
rect 506 958 522 1000
rect 562 958 574 1000
rect 506 940 574 958
rect -720 824 1020 874
rect -328 696 -294 824
rect 566 698 600 824
rect -656 326 -594 342
rect -656 284 -642 326
rect -606 284 -594 326
rect -656 268 -594 284
rect 864 328 926 344
rect 864 286 878 328
rect 914 286 926 328
rect -484 238 756 272
rect 864 270 926 286
rect -718 44 -652 200
rect -484 188 -450 238
rect -292 194 -258 238
rect -100 190 -66 238
rect 126 148 160 238
rect 338 192 372 238
rect 530 194 564 238
rect 722 192 756 238
rect -598 -22 -564 52
rect 30 48 66 88
rect 222 48 256 86
rect 30 -22 256 48
rect 836 -22 870 54
rect 954 42 1020 198
rect -720 -74 1020 -22
rect -422 -166 -128 -150
rect -422 -234 -406 -166
rect -144 -234 -128 -166
rect -422 -252 -128 -234
rect 78 -170 206 -152
rect 78 -238 104 -170
rect 180 -238 206 -170
rect 78 -260 206 -238
rect 398 -164 696 -148
rect 398 -234 414 -164
rect 680 -234 696 -164
rect 398 -250 696 -234
<< viali >>
rect -286 958 -250 1000
rect 522 958 562 1000
rect -642 284 -640 326
rect -640 284 -606 326
rect 878 286 880 328
rect 880 286 914 328
rect -406 -168 -144 -166
rect -406 -234 -144 -168
rect 106 -238 180 -170
rect 414 -234 680 -164
<< metal1 >>
rect -302 1000 -234 1016
rect -302 958 -286 1000
rect -250 958 -234 1000
rect -302 940 -234 958
rect 506 1000 574 1016
rect 506 958 522 1000
rect 562 958 574 1000
rect 506 940 574 958
rect -656 326 -594 342
rect -248 326 -200 592
rect 472 326 520 620
rect 864 328 926 344
rect 864 326 878 328
rect -718 284 -642 326
rect -606 284 -160 326
rect -656 268 -594 284
rect -692 190 -648 212
rect -390 154 -352 284
rect -198 150 -160 284
rect 434 286 878 326
rect 914 326 926 328
rect 914 286 1020 326
rect 434 284 1020 286
rect 434 188 470 284
rect 624 192 660 284
rect 864 270 926 284
rect -422 -166 -128 -150
rect -422 -234 -406 -166
rect -144 -234 -128 -166
rect -422 -254 -128 -234
rect 78 -170 206 -152
rect 78 -238 106 -170
rect 180 -238 206 -170
rect 78 -258 206 -238
rect 398 -164 696 -148
rect 398 -234 414 -164
rect 680 -234 696 -164
rect 398 -250 696 -234
use sky130_fd_pr__nfet_01v8_8FHE5N  sky130_fd_pr__nfet_01v8_8FHE5N_0
timestamp 1646423143
transform 1 0 143 0 1 126
box -125 -76 125 76
use sky130_fd_pr__nfet_01v8_F5U58G#1  sky130_fd_pr__nfet_01v8_F5U58G_0
timestamp 1646431323
transform 1 0 -625 0 1 116
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_F5U58G#1  sky130_fd_pr__nfet_01v8_F5U58G_1
timestamp 1646431323
transform 1 0 897 0 1 120
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_G6PLX8  sky130_fd_pr__nfet_01v8_G6PLX8_0
timestamp 1646422066
transform 1 0 -275 0 1 122
box -221 -126 221 150
use sky130_fd_pr__nfet_01v8_G6PLX8  sky130_fd_pr__nfet_01v8_G6PLX8_1
timestamp 1646422066
transform 1 0 547 0 1 122
box -221 -126 221 150
use sky130_fd_pr__pfet_01v8_RFM3CD#0  sky130_fd_pr__pfet_01v8_RFM3CD_0
timestamp 1646431323
transform 1 0 -267 0 1 648
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_RFM3CD#0  sky130_fd_pr__pfet_01v8_RFM3CD_1
timestamp 1646431323
transform 1 0 539 0 1 648
box -109 -162 109 162
<< end >>
