magic
tech sky130A
magscale 1 2
timestamp 1646325283
<< nwell >>
rect 82 814 3088 860
rect 706 580 740 630
rect 898 580 932 626
rect 1090 580 1124 630
rect 1282 580 1316 626
rect 1474 580 1508 628
rect 1666 580 1700 626
rect 598 546 1858 580
<< poly >>
rect 82 816 3088 862
rect 468 490 596 574
rect 468 436 498 490
rect 560 436 596 490
rect 468 358 596 436
<< polycont >>
rect 498 436 560 490
<< locali >>
rect -14 902 3188 954
rect 32 770 70 902
rect 224 770 262 902
rect 416 770 454 902
rect 608 768 646 902
rect 800 766 838 902
rect 992 768 1030 902
rect 1186 770 1224 902
rect 1376 766 1414 902
rect 1568 768 1606 902
rect 1760 766 1798 902
rect 1954 768 1992 902
rect 2146 768 2184 902
rect 2336 766 2374 902
rect 2528 760 2566 902
rect 2720 766 2758 902
rect 2912 768 2950 902
rect 3104 768 3142 902
rect 130 580 164 628
rect 322 580 356 630
rect 514 580 548 626
rect 706 580 740 630
rect 898 580 932 626
rect 1090 580 1124 630
rect 1282 580 1316 626
rect 1474 580 1508 628
rect 1666 580 1700 626
rect 1858 580 1892 628
rect 2050 580 2084 632
rect 128 546 2084 580
rect 2050 494 2084 546
rect 1944 492 2084 494
rect 2242 492 2276 634
rect 2434 492 2468 632
rect 2626 492 2660 630
rect 2818 492 2852 628
rect 3010 492 3044 632
rect -14 436 498 490
rect 560 436 576 490
rect 1944 436 3188 492
rect -14 434 152 436
rect 1944 390 2062 436
rect 512 354 2062 390
rect 514 314 552 354
rect 706 300 744 354
rect 900 304 938 354
rect 1090 302 1128 354
rect 1282 308 1320 354
rect 1476 304 1514 354
rect 1666 308 1704 354
rect 1858 308 1896 354
rect -14 0 3188 52
use sky130_fd_pr__nfet_01v8_VJWT33  sky130_fd_pr__nfet_01v8_VJWT33_0
timestamp 1646295505
transform 1 0 1205 0 1 242
box -797 -218 797 138
use sky130_fd_pr__pfet_01v8_3M44SC  sky130_fd_pr__pfet_01v8_3M44SC_0
timestamp 1646261959
transform 1 0 1587 0 1 700
box -1601 -200 1601 200
<< end >>
