magic
tech sky130A
magscale 1 2
timestamp 1646259600
<< error_p >>
rect -353 262 449 300
rect -449 -262 449 262
rect -449 -300 353 -262
<< nwell >>
rect -353 262 449 300
rect -449 -262 449 262
rect -449 -300 353 -262
<< pmos >>
rect -351 -200 -321 200
rect -255 -200 -225 200
rect -159 -200 -129 200
rect -63 -200 -33 200
rect 33 -200 63 200
rect 129 -200 159 200
rect 225 -200 255 200
rect 321 -200 351 200
<< pdiff >>
rect -409 144 -351 200
rect -413 132 -351 144
rect -413 -132 -401 132
rect -367 -132 -351 132
rect -413 -144 -351 -132
rect -409 -200 -351 -144
rect -321 132 -255 200
rect -321 -132 -305 132
rect -271 -132 -255 132
rect -321 -200 -255 -132
rect -225 132 -159 200
rect -225 -132 -209 132
rect -175 -132 -159 132
rect -225 -200 -159 -132
rect -129 132 -63 200
rect -129 -132 -113 132
rect -79 -132 -63 132
rect -129 -200 -63 -132
rect -33 132 33 200
rect -33 -132 -17 132
rect 17 -132 33 132
rect -33 -200 33 -132
rect 63 132 129 200
rect 63 -132 79 132
rect 113 -132 129 132
rect 63 -200 129 -132
rect 159 132 225 200
rect 159 -132 175 132
rect 209 -132 225 132
rect 159 -200 225 -132
rect 255 132 321 200
rect 255 -132 271 132
rect 305 -132 321 132
rect 255 -200 321 -132
rect 351 144 409 200
rect 351 132 413 144
rect 351 -132 367 132
rect 401 -132 413 132
rect 351 -144 413 -132
rect 351 -200 409 -144
<< pdiffc >>
rect -401 -132 -367 132
rect -305 -132 -271 132
rect -209 -132 -175 132
rect -113 -132 -79 132
rect -17 -132 17 132
rect 79 -132 113 132
rect 175 -132 209 132
rect 271 -132 305 132
rect 367 -132 401 132
<< poly >>
rect -273 281 -207 297
rect -273 247 -257 281
rect -223 247 -207 281
rect -273 231 -207 247
rect -81 281 -15 297
rect -81 247 -65 281
rect -31 247 -15 281
rect -81 231 -15 247
rect 111 281 177 297
rect 111 247 127 281
rect 161 247 177 281
rect 111 231 177 247
rect 303 281 369 297
rect 303 247 319 281
rect 353 247 369 281
rect 303 231 369 247
rect -351 200 -321 226
rect -255 200 -225 231
rect -159 200 -129 226
rect -63 200 -33 231
rect 33 200 63 226
rect 129 200 159 231
rect 225 200 255 226
rect 321 200 351 231
rect -351 -231 -321 -200
rect -255 -226 -225 -200
rect -159 -231 -129 -200
rect -63 -226 -33 -200
rect 33 -231 63 -200
rect 129 -226 159 -200
rect 225 -231 255 -200
rect 321 -226 351 -200
rect -369 -247 -303 -231
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -369 -297 -303 -281
rect -177 -247 -111 -231
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect -177 -297 -111 -281
rect 15 -247 81 -231
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 15 -297 81 -281
rect 207 -247 273 -231
rect 207 -281 223 -247
rect 257 -281 273 -247
rect 207 -297 273 -281
<< polycont >>
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
<< locali >>
rect -273 247 -257 281
rect -223 247 -207 281
rect -81 247 -65 281
rect -31 247 -15 281
rect 111 247 127 281
rect 161 247 177 281
rect 303 247 319 281
rect 353 247 369 281
rect -401 132 -367 148
rect -401 -148 -367 -132
rect -305 132 -271 148
rect -305 -148 -271 -132
rect -209 132 -175 148
rect -209 -148 -175 -132
rect -113 132 -79 148
rect -113 -148 -79 -132
rect -17 132 17 148
rect -17 -148 17 -132
rect 79 132 113 148
rect 79 -148 113 -132
rect 175 132 209 148
rect 175 -148 209 -132
rect 271 132 305 148
rect 271 -148 305 -132
rect 367 132 401 148
rect 367 -148 401 -132
rect -369 -281 -353 -247
rect -319 -281 -303 -247
rect -177 -281 -161 -247
rect -127 -281 -111 -247
rect 15 -281 31 -247
rect 65 -281 81 -247
rect 207 -281 223 -247
rect 257 -281 273 -247
<< viali >>
rect -257 247 -223 281
rect -65 247 -31 281
rect 127 247 161 281
rect 319 247 353 281
rect -401 -132 -367 132
rect -305 -132 -271 132
rect -209 -132 -175 132
rect -113 -132 -79 132
rect -17 -132 17 132
rect 79 -132 113 132
rect 175 -132 209 132
rect 271 -132 305 132
rect 367 -132 401 132
rect -353 -281 -319 -247
rect -161 -281 -127 -247
rect 31 -281 65 -247
rect 223 -281 257 -247
<< metal1 >>
rect -269 281 -211 287
rect -269 247 -257 281
rect -223 247 -211 281
rect -269 241 -211 247
rect -77 281 -19 287
rect -77 247 -65 281
rect -31 247 -19 281
rect -77 241 -19 247
rect 115 281 173 287
rect 115 247 127 281
rect 161 247 173 281
rect 115 241 173 247
rect 307 281 365 287
rect 307 247 319 281
rect 353 247 365 281
rect 307 241 365 247
rect -407 132 -361 144
rect -407 -132 -401 132
rect -367 -132 -361 132
rect -407 -144 -361 -132
rect -311 132 -265 144
rect -311 -132 -305 132
rect -271 -132 -265 132
rect -311 -144 -265 -132
rect -215 132 -169 144
rect -215 -132 -209 132
rect -175 -132 -169 132
rect -215 -144 -169 -132
rect -119 132 -73 144
rect -119 -132 -113 132
rect -79 -132 -73 132
rect -119 -144 -73 -132
rect -23 132 23 144
rect -23 -132 -17 132
rect 17 -132 23 132
rect -23 -144 23 -132
rect 73 132 119 144
rect 73 -132 79 132
rect 113 -132 119 132
rect 73 -144 119 -132
rect 169 132 215 144
rect 169 -132 175 132
rect 209 -132 215 132
rect 169 -144 215 -132
rect 265 132 311 144
rect 265 -132 271 132
rect 305 -132 311 132
rect 265 -144 311 -132
rect 361 132 407 144
rect 361 -132 367 132
rect 401 -132 407 132
rect 361 -144 407 -132
rect -365 -247 -307 -241
rect -365 -281 -353 -247
rect -319 -281 -307 -247
rect -365 -287 -307 -281
rect -173 -247 -115 -241
rect -173 -281 -161 -247
rect -127 -281 -115 -247
rect -173 -287 -115 -281
rect 19 -247 77 -241
rect 19 -281 31 -247
rect 65 -281 77 -247
rect 19 -287 77 -281
rect 211 -247 269 -241
rect 211 -281 223 -247
rect 257 -281 269 -247
rect 211 -287 269 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.15 m 1 nf 8 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
