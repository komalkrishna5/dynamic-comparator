magic
tech sky130A
timestamp 1645025748
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 2 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 20 viadrn 20 viagate 20 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
