magic
tech sky130A
magscale 1 2
timestamp 1646423143
<< nmos >>
rect -63 -50 -33 50
rect 33 -50 63 50
<< ndiff >>
rect -121 39 -63 50
rect -125 27 -63 39
rect -125 -27 -113 27
rect -79 -27 -63 27
rect -125 -39 -63 -27
rect -121 -50 -63 -39
rect -33 27 33 50
rect -33 -27 -17 27
rect 17 -27 33 27
rect -33 -50 33 -27
rect 63 39 121 50
rect 63 27 125 39
rect 63 -27 79 27
rect 113 -27 125 27
rect 63 -39 125 -27
rect 63 -50 121 -39
<< ndiffc >>
rect -113 -27 -79 27
rect -17 -27 17 27
rect 79 -27 113 27
<< poly >>
rect -63 50 -33 76
rect 33 50 63 76
rect -63 -76 -33 -50
rect 33 -76 63 -50
<< locali >>
rect -113 27 -79 43
rect -113 -43 -79 -27
rect -17 27 17 43
rect -17 -43 17 -27
rect 79 27 113 43
rect 79 -43 113 -27
<< viali >>
rect -113 -27 -79 27
rect -17 -27 17 27
rect 79 -27 113 27
<< metal1 >>
rect -119 27 -73 39
rect -119 -27 -113 27
rect -79 -27 -73 27
rect -119 -39 -73 -27
rect -23 27 23 39
rect -23 -27 -17 27
rect 17 -27 23 27
rect -23 -39 23 -27
rect 73 27 119 39
rect 73 -27 79 27
rect 113 -27 119 27
rect 73 -39 119 -27
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.150 m 1 nf 2 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
