magic
tech sky130A
magscale 1 2
timestamp 1647011741
<< nwell >>
rect 782 5052 940 5336
rect -348 3152 148 3568
rect 178 2078 1624 2402
rect 176 778 406 1044
<< psubdiff >>
rect 86 128 158 152
rect 86 -24 158 0
<< nsubdiff >>
rect 810 5270 888 5294
rect 810 5066 888 5090
rect -42 3424 26 3448
rect -42 3276 26 3300
rect 332 2308 416 2332
rect 332 2138 416 2162
rect 194 1008 312 1032
rect 194 784 312 808
<< psubdiffcont >>
rect 86 0 158 128
<< nsubdiffcont >>
rect 810 5090 888 5270
rect -42 3300 26 3424
rect 332 2162 416 2308
rect 194 808 312 1008
<< poly >>
rect 154 4922 262 4948
rect 154 4870 178 4922
rect 228 4916 262 4922
rect 228 4872 682 4916
rect 228 4870 262 4872
rect 154 4842 262 4870
rect 652 4812 682 4872
rect 1368 4580 1442 4600
rect 1368 4578 1384 4580
rect 1048 4532 1384 4578
rect 1426 4532 1442 4580
rect 1368 4518 1442 4532
rect 2540 4450 2636 4468
rect 2540 4406 2576 4450
rect 2618 4406 2636 4450
rect 2540 4382 2636 4406
rect 760 3868 984 3890
rect 760 3798 828 3868
rect 928 3798 984 3868
rect 760 3478 984 3798
rect 510 2556 584 2576
rect 510 2518 530 2556
rect 566 2518 584 2556
rect 510 2494 584 2518
rect 1090 2556 1164 2576
rect 1090 2518 1110 2556
rect 1146 2518 1164 2556
rect 1090 2494 1164 2518
rect 530 2348 560 2494
rect 1112 2350 1142 2494
rect 818 1490 848 1606
rect 816 1322 848 1490
rect 814 1276 850 1322
rect 802 1260 870 1276
rect 802 1218 818 1260
rect 858 1218 870 1260
rect 802 1200 870 1218
<< polycont >>
rect 178 4870 228 4922
rect 1384 4532 1426 4580
rect 2576 4406 2618 4450
rect 828 3798 928 3868
rect 530 2518 566 2556
rect 1110 2518 1146 2556
rect 818 1218 858 1260
<< locali >>
rect 3694 6986 4172 7104
rect 3694 6924 3812 6986
rect 3692 6790 3812 6924
rect 3694 6736 3812 6790
rect 4076 6736 4172 6986
rect 3694 6626 4172 6736
rect 3694 6230 4172 6348
rect 3694 6168 3812 6230
rect 2514 6034 3812 6168
rect 3694 5980 3812 6034
rect 4076 5980 4172 6230
rect 3694 5870 4172 5980
rect -2594 5556 -1352 5562
rect -2594 5526 -1346 5556
rect -2592 4638 -1346 5526
rect 3336 5454 4532 5556
rect 3336 5414 3428 5454
rect 3334 5410 3428 5414
rect 2612 5408 3428 5410
rect 396 5398 3428 5408
rect 822 5286 880 5374
rect 1148 5352 3428 5398
rect 810 5270 888 5286
rect 810 5074 888 5090
rect 3336 5214 3428 5352
rect 3652 5214 4228 5454
rect 4452 5214 4532 5454
rect 154 4922 262 4948
rect 154 4870 178 4922
rect 228 4870 262 4922
rect 154 4840 262 4870
rect 514 4852 776 4920
rect 1090 4862 1190 4936
rect 3336 4908 4532 5214
rect 2658 4858 4532 4908
rect -2592 4292 -2512 4638
rect -2262 4292 -1712 4638
rect -1462 4508 -1346 4638
rect 1368 4580 1442 4600
rect 1368 4532 1384 4580
rect 1426 4532 1442 4580
rect 1368 4518 1442 4532
rect -1462 4454 424 4508
rect -1462 4292 -1346 4454
rect 2178 4438 2308 4462
rect 2178 4362 2202 4438
rect 2274 4362 2308 4438
rect 2462 4456 2638 4470
rect 2462 4446 2568 4456
rect 2462 4400 2480 4446
rect 2530 4400 2568 4446
rect 2624 4400 2638 4456
rect 2462 4382 2638 4400
rect 2178 4336 2308 4362
rect -2592 4010 -1346 4292
rect -2592 3956 2294 4010
rect -2592 2826 -1346 3956
rect 798 3868 954 3892
rect 798 3798 828 3868
rect 928 3798 954 3868
rect 798 3778 954 3798
rect -50 3698 32 3710
rect -50 3638 -38 3698
rect 20 3638 32 3698
rect -50 3622 32 3638
rect 3336 3696 4532 4858
rect -28 3440 10 3622
rect 3336 3456 3428 3696
rect 3652 3456 4228 3696
rect 4452 3456 4532 3696
rect -42 3424 26 3440
rect -42 3284 26 3300
rect 1646 3028 1702 3128
rect 1646 2994 1656 3028
rect 1692 2994 1702 3028
rect 1646 2992 1702 2994
rect 2318 2848 2670 2898
rect 2318 2844 2386 2848
rect -2592 2480 -2512 2826
rect -2262 2480 -1712 2826
rect -1462 2764 -1346 2826
rect 2320 2772 2386 2844
rect -1462 2762 -34 2764
rect -1462 2710 84 2762
rect 2318 2716 2386 2772
rect -1462 2480 -1346 2710
rect -32 2688 84 2710
rect -32 2636 146 2688
rect -32 2634 84 2636
rect -882 2540 -530 2590
rect 2320 2586 2386 2716
rect 2612 2772 2670 2848
rect 2612 2716 2674 2772
rect 2612 2586 2670 2716
rect -882 2536 -814 2540
rect -2592 1726 -1346 2480
rect -880 2278 -814 2536
rect -588 2278 -530 2540
rect 512 2556 582 2572
rect 512 2518 530 2556
rect 566 2518 582 2556
rect 512 2502 582 2518
rect 1092 2556 1162 2572
rect 1092 2518 1110 2556
rect 1146 2518 1162 2556
rect 2320 2536 2670 2586
rect 3336 2536 4532 3456
rect 1092 2502 1162 2518
rect 3336 2464 3428 2536
rect 80 2410 280 2464
rect 1382 2462 2058 2464
rect 3282 2462 3428 2464
rect 1382 2408 3428 2462
rect 2098 2406 3276 2408
rect -880 2228 -530 2278
rect 332 2308 518 2334
rect 416 2162 518 2308
rect 332 2136 518 2162
rect 3336 2296 3428 2408
rect 3652 2296 4228 2536
rect 4452 2296 4532 2536
rect -2592 1380 -2512 1726
rect -2262 1380 -1712 1726
rect -1462 1572 -1346 1726
rect -1462 1514 332 1572
rect 2320 1550 2670 1600
rect -1462 1380 -1346 1514
rect -2592 426 -1346 1380
rect -880 1358 -530 1408
rect -880 1096 -814 1358
rect -588 1096 -530 1358
rect 2320 1332 2386 1550
rect 2318 1288 2386 1332
rect 2612 1288 2670 1550
rect 802 1260 870 1276
rect 2318 1274 2670 1288
rect 802 1218 818 1260
rect 858 1218 870 1260
rect 2320 1238 2670 1274
rect 802 1200 870 1218
rect 3336 1236 4532 2296
rect 3336 1140 3428 1236
rect 1650 1138 2318 1140
rect 2670 1138 3428 1140
rect -880 1046 -530 1096
rect -270 1084 62 1134
rect 1650 1082 3428 1138
rect 194 1008 426 1024
rect 312 830 426 1008
rect 3336 996 3428 1082
rect 3652 996 4228 1236
rect 4452 996 4532 1236
rect 194 792 312 808
rect -2592 80 -2512 426
rect -2262 80 -1712 426
rect -1462 238 -1346 426
rect -1462 186 26 238
rect 120 202 158 230
rect -1462 80 -1346 186
rect -2592 -824 -1346 80
rect 86 128 158 202
rect 86 -16 158 0
rect -880 -102 -530 -52
rect -880 -364 -814 -102
rect -588 -150 -530 -102
rect -588 -364 -530 -322
rect -880 -416 -530 -364
rect 3336 -788 4532 996
<< viali >>
rect -154 6788 -118 6894
rect 780 6778 816 6882
rect 1610 6784 1644 6886
rect 2252 6784 2288 6886
rect 3812 6736 4076 6986
rect 96 6058 130 6160
rect 1028 6060 1062 6162
rect 1802 6060 1836 6162
rect 3812 5980 4076 6230
rect 3428 5214 3652 5454
rect 4228 5214 4452 5454
rect 178 4870 228 4922
rect -2512 4292 -2262 4638
rect -1712 4292 -1462 4638
rect 1384 4532 1426 4580
rect 2202 4362 2274 4438
rect 2568 4450 2624 4456
rect 2480 4400 2530 4446
rect 2568 4406 2576 4450
rect 2576 4406 2618 4450
rect 2618 4406 2624 4450
rect 2568 4400 2624 4406
rect 828 3798 928 3868
rect -38 3638 20 3698
rect 3428 3456 3652 3696
rect 4228 3456 4452 3696
rect 306 3078 356 3124
rect 1384 3078 1434 3124
rect 1656 2994 1692 3028
rect -2512 2480 -2262 2826
rect -1712 2480 -1462 2826
rect 2386 2586 2612 2848
rect -814 2278 -588 2540
rect 530 2518 566 2556
rect 1110 2518 1146 2556
rect 3428 2296 3652 2536
rect 4228 2296 4452 2536
rect -2512 1380 -2262 1726
rect -1712 1380 -1462 1726
rect -814 1096 -588 1358
rect 2386 1288 2612 1550
rect 818 1218 858 1260
rect 3428 996 3652 1236
rect 4228 996 4452 1236
rect -2512 80 -2262 426
rect -1712 80 -1462 426
rect -814 -364 -588 -102
<< metal1 >>
rect -2282 6952 -1768 7064
rect -2282 6686 -2174 6952
rect -1874 6916 -1768 6952
rect 3692 6986 4174 7106
rect -1318 6916 -104 6920
rect -1874 6894 -104 6916
rect -1874 6788 -154 6894
rect -118 6788 -104 6894
rect -1874 6766 -104 6788
rect -64 6882 822 6904
rect -64 6778 780 6882
rect 816 6778 822 6882
rect -64 6766 822 6778
rect -1874 6762 -590 6766
rect 88 6764 822 6766
rect 876 6886 1666 6904
rect 876 6784 1610 6886
rect 1644 6784 1666 6886
rect 876 6764 1666 6784
rect 1702 6886 2310 6902
rect 3692 6896 3812 6986
rect 1702 6784 2252 6886
rect 2288 6784 2310 6886
rect 1702 6770 2310 6784
rect 2350 6764 3812 6896
rect 3202 6762 3812 6764
rect -1874 6686 -1768 6762
rect -2282 6560 -1768 6686
rect 3692 6736 3812 6762
rect 4076 6736 4174 6986
rect 3692 6624 4174 6736
rect -2282 6226 -1768 6338
rect -2282 5960 -2174 6226
rect -1874 6172 -1768 6226
rect 3692 6230 4174 6350
rect -1874 6168 -614 6172
rect -1874 6050 34 6168
rect 84 6160 968 6168
rect 84 6058 96 6160
rect 130 6058 968 6160
rect 84 6050 968 6058
rect 1012 6162 1740 6174
rect 1012 6060 1028 6162
rect 1062 6060 1740 6162
rect 1012 6054 1740 6060
rect 1790 6162 2452 6178
rect 1790 6060 1802 6162
rect 1836 6060 2452 6162
rect -1874 6046 -614 6050
rect 1790 6046 2452 6060
rect -1874 5960 -1768 6046
rect -2282 5834 -1768 5960
rect 3692 5980 3812 6230
rect 4076 5980 4174 6230
rect 3692 5868 4174 5980
rect 3358 5454 3714 5514
rect 3358 5214 3428 5454
rect 3652 5214 3714 5454
rect 3358 5148 3714 5214
rect 4156 5454 4514 5514
rect 4156 5214 4228 5454
rect 4452 5214 4514 5454
rect 4156 5148 4514 5214
rect 154 4938 262 4948
rect -210 4922 262 4938
rect -210 4870 178 4922
rect 228 4870 262 4922
rect -210 4854 262 4870
rect -210 4776 -126 4854
rect 154 4840 262 4854
rect -2570 4638 -2204 4684
rect -2570 4292 -2512 4638
rect -2262 4292 -2204 4638
rect -2570 4226 -2204 4292
rect -1770 4638 -1404 4684
rect -208 4680 -128 4776
rect -1770 4292 -1712 4638
rect -1462 4292 -1404 4638
rect -1770 4226 -1404 4292
rect -210 3792 -128 4680
rect 1368 4580 1442 4600
rect 1368 4532 1384 4580
rect 1426 4570 1972 4580
rect 1426 4534 1976 4570
rect 1426 4532 1442 4534
rect 1368 4518 1442 4532
rect 1886 4488 1976 4534
rect 1890 3922 1972 4488
rect 2538 4468 2638 4470
rect 2178 4438 2308 4462
rect 2178 4362 2202 4438
rect 2274 4362 2308 4438
rect 2462 4456 2638 4468
rect 2462 4400 2480 4456
rect 2536 4400 2568 4456
rect 2624 4400 2638 4456
rect 2462 4382 2638 4400
rect 2178 4336 2308 4362
rect -208 3128 -128 3792
rect 798 3868 954 3892
rect 798 3798 828 3868
rect 928 3798 954 3868
rect 798 3778 954 3798
rect -50 3698 32 3710
rect 804 3702 1042 3728
rect 804 3698 866 3702
rect -50 3638 -38 3698
rect 20 3638 866 3698
rect -50 3636 866 3638
rect -50 3622 32 3636
rect 804 3622 866 3636
rect 970 3622 1042 3702
rect 804 3600 1042 3622
rect 272 3128 374 3144
rect -208 3124 374 3128
rect -208 3078 306 3124
rect 356 3078 374 3124
rect -208 3072 374 3078
rect -2570 2826 -2204 2876
rect -2570 2480 -2512 2826
rect -2262 2480 -2204 2826
rect -2570 2414 -2204 2480
rect -1770 2826 -1404 2876
rect -1770 2480 -1712 2826
rect -1462 2480 -1404 2826
rect -1770 2414 -1404 2480
rect -882 2540 -530 2590
rect -882 2278 -814 2540
rect -588 2278 -530 2540
rect -882 2228 -530 2278
rect -2570 1726 -2204 1776
rect -2570 1380 -2512 1726
rect -2262 1380 -2204 1726
rect -2570 1314 -2204 1380
rect -1770 1726 -1404 1776
rect -1770 1380 -1712 1726
rect -1462 1380 -1404 1726
rect -1770 1314 -1404 1380
rect -882 1358 -530 1408
rect -882 1096 -814 1358
rect -588 1096 -530 1358
rect -882 1046 -530 1096
rect -2570 426 -2204 476
rect -2570 80 -2512 426
rect -2262 80 -2204 426
rect -2570 14 -2204 80
rect -1770 426 -1404 476
rect -1770 80 -1712 426
rect -1462 80 -1404 426
rect -208 398 -128 3072
rect 272 3030 374 3072
rect 1368 3124 1452 3144
rect 1368 3078 1384 3124
rect 1434 3122 1452 3124
rect 1892 3122 1972 3922
rect 3356 3696 3714 3756
rect 3356 3456 3428 3696
rect 3652 3456 3714 3696
rect 3356 3390 3714 3456
rect 4156 3696 4514 3756
rect 4156 3456 4228 3696
rect 4452 3456 4514 3696
rect 4156 3390 4514 3456
rect 1434 3078 1974 3122
rect 1368 3072 1974 3078
rect 1368 3060 1452 3072
rect 1646 3030 1704 3040
rect 272 3028 1704 3030
rect 272 2994 1656 3028
rect 1692 2994 1704 3028
rect 1892 3002 1974 3072
rect 272 2992 1704 2994
rect 1646 2980 1704 2992
rect 512 2564 582 2572
rect 512 2512 524 2564
rect 576 2512 582 2564
rect 512 2502 582 2512
rect 1092 2564 1162 2572
rect 1092 2512 1104 2564
rect 1156 2512 1162 2564
rect 1092 2502 1162 2512
rect -58 1930 306 1992
rect 1202 1938 1806 2000
rect -58 586 -2 1930
rect 260 1900 306 1930
rect 260 1888 304 1900
rect 802 1268 870 1276
rect 802 1210 810 1268
rect 866 1210 870 1268
rect 802 1200 870 1210
rect 1750 586 1806 1938
rect -58 544 40 586
rect 1716 544 1806 586
rect 1894 412 1974 3002
rect 2318 2848 2670 2898
rect 2318 2586 2386 2848
rect 2612 2586 2670 2848
rect 2318 2536 2670 2586
rect 3356 2536 3714 2596
rect 3356 2296 3428 2536
rect 3652 2296 3714 2536
rect 3356 2230 3714 2296
rect 4156 2536 4514 2596
rect 4156 2296 4228 2536
rect 4452 2296 4514 2536
rect 4156 2230 4514 2296
rect 2318 1550 2670 1600
rect 2318 1288 2386 1550
rect 2612 1288 2670 1550
rect 2318 1238 2670 1288
rect 3356 1236 3714 1298
rect 3356 996 3428 1236
rect 3652 996 3714 1236
rect 3356 930 3714 996
rect 4156 1236 4514 1298
rect 4156 996 4228 1236
rect 4452 996 4514 1236
rect 4156 930 4514 996
rect -208 342 70 398
rect 1638 356 1974 412
rect -1770 14 -1404 80
rect -882 -102 -530 -52
rect -882 -364 -814 -102
rect -588 -364 -530 -102
rect 296 -116 590 108
rect 1116 -116 1416 112
rect -882 -416 -530 -364
<< via1 >>
rect -2174 6686 -1874 6952
rect 3812 6736 4076 6986
rect -2174 5960 -1874 6226
rect 3812 5980 4076 6230
rect 3428 5214 3652 5454
rect 4228 5214 4452 5454
rect -2512 4292 -2262 4638
rect -1712 4292 -1462 4638
rect 2202 4362 2274 4438
rect 2480 4446 2536 4456
rect 2480 4400 2530 4446
rect 2530 4400 2536 4446
rect 2568 4400 2624 4456
rect 828 3798 928 3868
rect 866 3622 970 3702
rect -2512 2480 -2262 2826
rect -1712 2480 -1462 2826
rect -814 2278 -588 2540
rect -2512 1380 -2262 1726
rect -1712 1380 -1462 1726
rect -814 1096 -588 1358
rect -2512 80 -2262 426
rect -1712 80 -1462 426
rect 3428 3456 3652 3696
rect 4228 3456 4452 3696
rect 524 2556 576 2564
rect 524 2518 530 2556
rect 530 2518 566 2556
rect 566 2518 576 2556
rect 524 2512 576 2518
rect 1104 2556 1156 2564
rect 1104 2518 1110 2556
rect 1110 2518 1146 2556
rect 1146 2518 1156 2556
rect 1104 2512 1156 2518
rect 424 1206 480 1268
rect 810 1260 866 1268
rect 810 1218 818 1260
rect 818 1218 858 1260
rect 858 1218 866 1260
rect 810 1210 866 1218
rect 1234 1210 1290 1268
rect 2386 2586 2612 2848
rect 3428 2296 3652 2536
rect 4228 2296 4452 2536
rect 2386 1318 2612 1550
rect 2386 1288 2610 1318
rect 3428 996 3652 1236
rect 4228 996 4452 1236
rect -814 -364 -588 -102
rect 812 10 910 98
<< metal2 >>
rect -2282 6952 -1768 7064
rect -2282 6686 -2174 6952
rect -1874 6686 -1768 6952
rect -2282 6560 -1768 6686
rect 3692 6986 4174 7106
rect 3692 6736 3812 6986
rect 4076 6736 4174 6986
rect 3692 6624 4174 6736
rect -2282 6226 -1768 6338
rect -2282 5960 -2174 6226
rect -1874 5960 -1768 6226
rect -2282 5834 -1768 5960
rect 3692 6230 4174 6350
rect 3692 5980 3812 6230
rect 4076 5980 4174 6230
rect 3692 5868 4174 5980
rect 3328 5454 4532 5558
rect 3328 5214 3428 5454
rect 3652 5214 4228 5454
rect 4452 5214 4532 5454
rect -2570 4638 -2204 4684
rect -2570 4292 -2512 4638
rect -2262 4292 -2204 4638
rect -2570 4226 -2204 4292
rect -1770 4638 -1404 4684
rect -1770 4292 -1712 4638
rect -1462 4292 -1404 4638
rect 2538 4468 2638 4470
rect -1770 4226 -1404 4292
rect 798 4438 2308 4462
rect 798 4362 2202 4438
rect 2274 4362 2308 4438
rect 2462 4456 2638 4468
rect 2462 4400 2480 4456
rect 2536 4400 2568 4456
rect 2624 4400 2638 4456
rect 2462 4382 2638 4400
rect 798 4336 2308 4362
rect 798 3868 956 4336
rect 798 3798 828 3868
rect 928 3798 956 3868
rect 798 3778 956 3798
rect 804 3702 1032 3718
rect 804 3622 866 3702
rect 970 3686 1032 3702
rect 3328 3696 4532 5214
rect 3328 3686 3428 3696
rect 970 3622 3428 3686
rect 804 3620 3428 3622
rect 804 3602 1032 3620
rect 3328 3456 3428 3620
rect 3652 3456 4228 3696
rect 4452 3456 4532 3696
rect -2570 2826 -2204 2876
rect -2570 2480 -2512 2826
rect -2262 2480 -2204 2826
rect -2570 2414 -2204 2480
rect -1770 2826 -1404 2876
rect -1770 2480 -1712 2826
rect -1462 2480 -1404 2826
rect -1770 2414 -1404 2480
rect -920 2558 -518 2942
rect 2278 2848 2680 2944
rect 2278 2586 2386 2848
rect 2612 2586 2680 2848
rect 2278 2580 2680 2586
rect 1156 2578 2680 2580
rect 510 2564 584 2576
rect 510 2558 524 2564
rect -920 2540 524 2558
rect -920 2278 -814 2540
rect -588 2512 524 2540
rect 576 2512 584 2564
rect -588 2510 584 2512
rect -588 2278 -518 2510
rect 510 2494 584 2510
rect 1090 2564 2680 2578
rect 1090 2512 1104 2564
rect 1156 2526 2680 2564
rect 1156 2512 1164 2526
rect 1090 2494 1164 2512
rect -920 2092 -518 2278
rect 2278 2096 2680 2526
rect -920 2026 370 2092
rect -2570 1726 -2204 1776
rect -2570 1380 -2512 1726
rect -2262 1380 -2204 1726
rect -2570 1314 -2204 1380
rect -1770 1726 -1404 1776
rect -1770 1380 -1712 1726
rect -1462 1380 -1404 1726
rect -1770 1314 -1404 1380
rect -920 1358 -518 2026
rect 1320 2024 2680 2096
rect 2278 1550 2680 2024
rect 2278 1370 2386 1550
rect -920 1096 -814 1358
rect -588 1352 -518 1358
rect 800 1354 872 1356
rect 412 1352 872 1354
rect -588 1304 872 1352
rect -588 1096 -518 1304
rect 412 1268 486 1304
rect 412 1206 424 1268
rect 480 1206 486 1268
rect 412 1200 486 1206
rect 800 1268 872 1304
rect 1234 1320 2386 1370
rect 1234 1276 1294 1320
rect 800 1210 810 1268
rect 866 1210 872 1268
rect 800 1200 872 1210
rect 1226 1268 1294 1276
rect 1226 1210 1234 1268
rect 1290 1210 1294 1268
rect 1226 1200 1294 1210
rect 2278 1288 2386 1320
rect 2612 1318 2680 1550
rect 2610 1288 2680 1318
rect -2570 426 -2204 476
rect -2570 80 -2512 426
rect -2262 80 -2204 426
rect -2570 14 -2204 80
rect -1770 426 -1404 476
rect -1770 80 -1712 426
rect -1462 80 -1404 426
rect -1770 14 -1404 80
rect -920 -102 -518 1096
rect -920 -364 -814 -102
rect -588 -210 -518 -102
rect 794 98 928 110
rect 794 10 812 98
rect 910 10 928 98
rect 794 -210 928 10
rect -588 -300 930 -210
rect -588 -364 -518 -300
rect -920 -536 -518 -364
rect 2278 -536 2680 1288
rect 3328 2536 4532 3456
rect 3328 2296 3428 2536
rect 3652 2296 4228 2536
rect 4452 2296 4532 2536
rect 3328 1236 4532 2296
rect 3328 996 3428 1236
rect 3652 996 4228 1236
rect 4452 996 4532 1236
rect -920 -824 2682 -536
rect 3328 -788 4532 996
<< via2 >>
rect -2174 6686 -1874 6952
rect 3812 6736 4076 6986
rect -2174 5960 -1874 6226
rect 3812 5980 4076 6230
rect 3428 5214 3652 5454
rect 4228 5214 4452 5454
rect -2512 4292 -2262 4638
rect -1712 4292 -1462 4638
rect 2480 4400 2536 4456
rect 2568 4400 2624 4456
rect 3428 3456 3652 3696
rect 4228 3456 4452 3696
rect -2512 2480 -2262 2826
rect -1712 2480 -1462 2826
rect 2386 2586 2612 2848
rect -814 2278 -588 2540
rect -2512 1380 -2262 1726
rect -1712 1380 -1462 1726
rect -814 1096 -588 1358
rect 2386 1318 2612 1550
rect 2386 1288 2610 1318
rect -2512 80 -2262 426
rect -1712 80 -1462 426
rect -814 -364 -588 -102
rect 3428 2296 3652 2536
rect 4228 2296 4452 2536
rect 3428 996 3652 1236
rect 4228 996 4452 1236
<< metal3 >>
rect -2282 6952 -1768 7064
rect -2282 6686 -2174 6952
rect -1874 6686 -1768 6952
rect -2282 6560 -1768 6686
rect 3692 6986 4174 7106
rect 3692 6736 3812 6986
rect 4076 6736 4174 6986
rect 3692 6624 4174 6736
rect -2282 6226 -1768 6338
rect -2282 5960 -2174 6226
rect -1874 5960 -1768 6226
rect -2282 5834 -1768 5960
rect 3692 6230 4174 6350
rect 3692 5980 3812 6230
rect 4076 5980 4174 6230
rect 3692 5868 4174 5980
rect 3358 5454 3714 5514
rect 3358 5214 3428 5454
rect 3652 5214 3714 5454
rect 3358 5148 3714 5214
rect 4156 5454 4514 5514
rect 4156 5214 4228 5454
rect 4452 5214 4514 5454
rect 4156 5148 4514 5214
rect -2570 4638 -2204 4684
rect -2570 4292 -2512 4638
rect -2262 4292 -2204 4638
rect -2570 4226 -2204 4292
rect -1770 4638 -1404 4684
rect -1770 4292 -1712 4638
rect -1462 4292 -1404 4638
rect -1770 4226 -1404 4292
rect 2274 4456 2680 4584
rect 2274 4400 2480 4456
rect 2536 4400 2568 4456
rect 2624 4400 2680 4456
rect 2274 3802 2680 4400
rect 2274 3704 2684 3802
rect -2570 2826 -2204 2876
rect -2570 2480 -2512 2826
rect -2262 2480 -2204 2826
rect -2570 2414 -2204 2480
rect -1770 2826 -1404 2876
rect -1770 2480 -1712 2826
rect -1462 2480 -1404 2826
rect -1770 2414 -1404 2480
rect -924 2540 -510 2948
rect 2278 2944 2684 3704
rect 3356 3696 3714 3756
rect 3356 3456 3428 3696
rect 3652 3456 3714 3696
rect 3356 3390 3714 3456
rect 4156 3696 4514 3756
rect 4156 3456 4228 3696
rect 4452 3456 4514 3696
rect 4156 3390 4514 3456
rect -924 2278 -814 2540
rect -588 2278 -510 2540
rect -2570 1726 -2204 1776
rect -2570 1380 -2512 1726
rect -2262 1380 -2204 1726
rect -2570 1314 -2204 1380
rect -1770 1726 -1404 1776
rect -1770 1380 -1712 1726
rect -1462 1380 -1404 1726
rect -1770 1314 -1404 1380
rect -924 1358 -510 2278
rect -924 1096 -814 1358
rect -588 1096 -510 1358
rect -2570 426 -2204 476
rect -2570 80 -2512 426
rect -2262 80 -2204 426
rect -2570 14 -2204 80
rect -1770 426 -1404 476
rect -1770 80 -1712 426
rect -1462 80 -1404 426
rect -1770 14 -1404 80
rect -924 -102 -510 1096
rect -924 -364 -814 -102
rect -588 -364 -510 -102
rect -924 -556 -510 -364
rect 2276 2848 2684 2944
rect 2276 2586 2386 2848
rect 2612 2586 2684 2848
rect 2276 1550 2684 2586
rect 3356 2536 3714 2596
rect 3356 2296 3428 2536
rect 3652 2296 3714 2536
rect 3356 2230 3714 2296
rect 4156 2536 4514 2596
rect 4156 2296 4228 2536
rect 4452 2296 4514 2536
rect 4156 2230 4514 2296
rect 2276 1288 2386 1550
rect 2612 1318 2684 1550
rect 2610 1288 2684 1318
rect 2276 -110 2684 1288
rect 3356 1236 3714 1298
rect 3356 996 3428 1236
rect 3652 996 3714 1236
rect 3356 930 3714 996
rect 4156 1236 4514 1298
rect 4156 996 4228 1236
rect 4452 996 4514 1236
rect 4156 930 4514 996
rect 2276 -356 2682 -110
rect 2276 -556 2684 -356
rect -924 -646 2684 -556
rect -920 -824 2684 -646
<< via3 >>
rect -2174 6686 -1874 6952
rect 3812 6736 4076 6986
rect -2174 5960 -1874 6226
rect 3812 5980 4076 6230
rect 3428 5214 3652 5454
rect 4228 5214 4452 5454
rect -2512 4292 -2262 4638
rect -1712 4292 -1462 4638
rect -2512 2480 -2262 2826
rect -1712 2480 -1462 2826
rect 3428 3456 3652 3696
rect 4228 3456 4452 3696
rect -2512 1380 -2262 1726
rect -1712 1380 -1462 1726
rect -2512 80 -2262 426
rect -1712 80 -1462 426
rect 3428 2296 3652 2536
rect 4228 2296 4452 2536
rect 3428 996 3652 1236
rect 4228 996 4452 1236
<< metal4 >>
rect 3322 7412 4536 7550
rect 3322 7130 4538 7412
rect -2282 6952 -1768 7064
rect -2282 6686 -2174 6952
rect -1874 6686 -1768 6952
rect -2282 6560 -1768 6686
rect 3324 6986 4538 7130
rect 3324 6736 3812 6986
rect 4076 6736 4538 6986
rect -2282 6226 -1768 6338
rect -2282 5960 -2174 6226
rect -1874 5960 -1768 6226
rect -2282 5834 -1768 5960
rect 3324 6230 4538 6736
rect 3324 5980 3812 6230
rect 4076 5980 4538 6230
rect 3324 5454 4538 5980
rect 3324 5214 3428 5454
rect 3652 5214 4228 5454
rect 4452 5214 4538 5454
rect 3324 4778 4538 5214
rect -2570 4638 -2204 4684
rect -2570 4292 -2512 4638
rect -2262 4292 -2204 4638
rect -2570 4226 -2204 4292
rect -1770 4638 -1404 4684
rect -1770 4292 -1712 4638
rect -1462 4292 -1404 4638
rect -1770 4226 -1404 4292
rect 3336 3696 4532 4778
rect 3336 3456 3428 3696
rect 3652 3456 4228 3696
rect 4452 3456 4532 3696
rect -2570 2826 -2204 2876
rect -2570 2480 -2512 2826
rect -2262 2480 -2204 2826
rect -2570 2414 -2204 2480
rect -1770 2826 -1404 2876
rect -1770 2480 -1712 2826
rect -1462 2480 -1404 2826
rect -1770 2414 -1404 2480
rect 3336 2536 4532 3456
rect 3336 2296 3428 2536
rect 3652 2296 4228 2536
rect 4452 2296 4532 2536
rect -2570 1726 -2204 1776
rect -2570 1380 -2512 1726
rect -2262 1380 -2204 1726
rect -2570 1314 -2204 1380
rect -1770 1726 -1404 1776
rect -1770 1380 -1712 1726
rect -1462 1380 -1404 1726
rect -1770 1314 -1404 1380
rect 3336 1236 4532 2296
rect 3336 996 3428 1236
rect 3652 996 4228 1236
rect 4452 996 4532 1236
rect -2570 426 -2204 476
rect -2570 80 -2512 426
rect -2262 80 -2204 426
rect -2570 14 -2204 80
rect -1770 426 -1404 476
rect -1770 80 -1712 426
rect -1462 80 -1404 426
rect -1770 14 -1404 80
rect 3336 -788 4532 996
<< via4 >>
rect -2174 6686 -1874 6952
rect -2174 5960 -1874 6226
rect -2512 4292 -2262 4638
rect -1712 4292 -1462 4638
rect -2512 2480 -2262 2826
rect -1712 2480 -1462 2826
rect -2512 1380 -2262 1726
rect -1712 1380 -1462 1726
rect -2512 80 -2262 426
rect -1712 80 -1462 426
<< metal5 >>
rect -2612 7202 -1346 7550
rect -2612 7030 -1344 7202
rect -2592 6952 -1344 7030
rect -2592 6686 -2174 6952
rect -1874 6686 -1344 6952
rect -2592 6226 -1344 6686
rect -2592 5960 -2174 6226
rect -1874 5960 -1344 6226
rect -2592 5374 -1344 5960
rect -2592 4638 -1354 5374
rect -2592 4292 -2512 4638
rect -2262 4292 -1712 4638
rect -1462 4292 -1354 4638
rect -2592 2826 -1354 4292
rect -2592 2480 -2512 2826
rect -2262 2480 -1712 2826
rect -1462 2480 -1354 2826
rect -2592 1726 -1354 2480
rect -2592 1380 -2512 1726
rect -2262 1380 -1712 1726
rect -1462 1380 -1354 1726
rect -2592 426 -1354 1380
rect -2592 80 -2512 426
rect -2262 80 -1712 426
rect -1462 80 -1354 426
rect -2592 -824 -1354 80
use SR_latch  SR_latch_0 ~/mycomparator_copy1/layout/latch
timestamp 1646810677
transform 1 0 394 0 1 4454
box 0 0 872 948
use inv_W1  inv_W1_0 ~/mycomparator_copy1/layout/myinv_layout2
timestamp 1645263751
transform -1 0 2630 0 1 4030
box -100 -72 388 878
use latch_2  latch_2_0 ~/mycomparator/layout/latch
timestamp 1646831438
transform 1 0 86 0 1 2636
box 0 0 1602 1002
use preamp_part1  preamp_part1_0 ~/mycomparator/layout/preamp
timestamp 1646810354
transform 1 0 720 0 1 260
box -720 -260 1020 1016
use preamp_part2  preamp_part2_0 ~/mycomparator/layout/preamp
timestamp 1646810398
transform 1 0 138 0 1 1376
box 116 2 1282 1088
use sky130_fd_pr__diode_pw2nd_05v5_FT7GK8  sky130_fd_pr__diode_pw2nd_05v5_FT7GK8_0
timestamp 1646995406
transform 1 0 2400 0 1 6834
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT7GK8  sky130_fd_pr__diode_pw2nd_05v5_FT7GK8_1
timestamp 1646995406
transform 1 0 1758 0 1 6836
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT7GK8  sky130_fd_pr__diode_pw2nd_05v5_FT7GK8_2
timestamp 1646995406
transform 1 0 928 0 1 6830
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_FT7GK8  sky130_fd_pr__diode_pw2nd_05v5_FT7GK8_3
timestamp 1646995406
transform 1 0 -6 0 1 6840
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_KLAK3C  sky130_fd_pr__diode_pw2nd_05v5_KLAK3C_0
timestamp 1646995406
transform 1 0 2400 0 1 6112
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_KLAK3C  sky130_fd_pr__diode_pw2nd_05v5_KLAK3C_1
timestamp 1646995406
transform 1 0 1689 0 1 6111
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_KLAK3C  sky130_fd_pr__diode_pw2nd_05v5_KLAK3C_2
timestamp 1646995406
transform 1 0 915 0 1 6111
box -183 -183 183 183
use sky130_fd_pr__diode_pw2nd_05v5_KLAK3C  sky130_fd_pr__diode_pw2nd_05v5_KLAK3C_3
timestamp 1646995406
transform 1 0 -17 0 1 6109
box -183 -183 183 183
<< labels >>
rlabel metal1 440 -116 440 -116 5 Vn
rlabel metal1 1280 -116 1280 -116 5 Vp
rlabel locali 514 4862 514 4862 7 Outp
rlabel locali 1190 4896 1190 4896 3 Outn
rlabel metal3 990 -824 990 -824 5 CLK
rlabel metal5 -2092 -824 -2092 -824 5 GND
rlabel metal4 3792 -788 3792 -788 5 VDD
<< end >>
