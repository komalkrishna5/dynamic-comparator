magic
tech sky130A
magscale 1 2
timestamp 1645025748
<< error_p >>
rect 19 181 77 187
rect 19 147 31 181
rect 19 141 77 147
<< nwell >>
rect -317 -202 169 204
<< pmos >>
rect -63 -100 -33 100
rect 33 -100 63 100
<< pdiff >>
rect -139 62 -63 100
rect -139 -62 -113 62
rect -79 -62 -63 62
rect -139 -100 -63 -62
rect -33 62 33 100
rect -33 -62 -17 62
rect 17 -62 33 62
rect -33 -100 33 -62
rect 63 74 121 100
rect 63 62 125 74
rect 63 -62 79 62
rect 113 -62 125 62
rect 63 -74 125 -62
rect 63 -100 121 -74
<< pdiffc >>
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
<< nsubdiff >>
rect -267 100 -179 124
rect -179 -100 -139 100
rect -267 -124 -179 -100
<< nsubdiffcont >>
rect -267 -100 -179 100
<< poly >>
rect 15 181 81 197
rect 15 147 31 181
rect 65 147 81 181
rect 15 131 81 147
rect -63 100 -33 126
rect 33 100 63 131
rect -63 -130 -33 -100
rect 33 -126 63 -100
<< polycont >>
rect 31 147 65 181
<< locali >>
rect 15 147 31 181
rect 65 147 81 181
rect -267 100 -179 116
rect -113 62 -79 78
rect -113 -78 -79 -62
rect -17 62 17 78
rect -17 -78 17 -62
rect 79 62 113 78
rect 79 -78 113 -62
rect -267 -116 -179 -100
<< viali >>
rect 31 147 65 181
rect -113 -44 -79 44
rect -17 -44 17 44
rect 79 -44 113 44
<< metal1 >>
rect 19 181 77 187
rect 19 147 31 181
rect 65 147 77 181
rect 19 141 77 147
rect -119 44 -73 56
rect -119 -44 -113 44
rect -79 -44 -73 44
rect -119 -56 -73 -44
rect -23 44 23 56
rect -23 -44 -17 44
rect 17 -44 23 44
rect -23 -56 23 -44
rect 73 44 119 56
rect 73 -44 79 44
rect 113 -44 119 44
rect 73 -56 119 -44
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 2 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 50 viadrn 50 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
