magic
tech sky130A
magscale 1 2
timestamp 1646325197
<< nwell >>
rect 354 500 2050 954
<< poly >>
rect 466 816 1940 862
rect 848 498 892 584
rect 804 482 892 498
rect 804 446 820 482
rect 856 446 892 482
rect 804 430 892 446
rect 848 364 892 430
<< polycont >>
rect 820 446 856 482
<< locali >>
rect 354 902 2050 954
rect 416 770 454 902
rect 608 768 646 902
rect 800 766 838 902
rect 992 768 1030 902
rect 1186 770 1224 902
rect 1376 766 1414 902
rect 1568 768 1606 902
rect 1760 766 1798 902
rect 1954 768 1992 902
rect 514 580 548 626
rect 706 580 740 630
rect 898 580 932 626
rect 1090 580 1124 630
rect 1282 580 1316 626
rect 1474 580 1508 628
rect 1666 580 1700 626
rect 1858 580 1892 628
rect 512 546 1898 580
rect 1516 492 1664 546
rect 354 482 888 490
rect 354 446 820 482
rect 856 446 888 482
rect 354 436 888 446
rect 1516 436 2050 492
rect 1516 390 1668 436
rect 900 354 1668 390
rect 900 304 938 354
rect 1090 302 1128 354
rect 1282 308 1320 354
rect 1476 304 1514 354
rect 806 52 840 168
rect 998 52 1032 174
rect 1190 52 1224 168
rect 1382 52 1416 174
rect 1574 52 1608 170
rect 354 0 2050 52
use sky130_fd_pr__nfet_01v8_KZU588  sky130_fd_pr__nfet_01v8_KZU588_0
timestamp 1646318752
transform 1 0 1207 0 1 240
box -413 -162 413 150
use sky130_fd_pr__pfet_01v8_RL4NCG  sky130_fd_pr__pfet_01v8_RL4NCG_0
timestamp 1646319668
transform 1 0 1203 0 1 700
box -833 -200 833 200
<< end >>
