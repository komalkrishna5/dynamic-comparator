magic
tech sky130A
magscale 1 2
timestamp 1646318752
<< error_p >>
rect 321 134 351 150
rect 321 116 355 134
<< nmos >>
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
<< ndiff >>
rect -409 74 -351 100
rect -413 62 -351 74
rect -413 -62 -401 62
rect -367 -62 -351 62
rect -413 -74 -351 -62
rect -409 -100 -351 -74
rect -321 62 -255 100
rect -321 -62 -305 62
rect -271 -62 -255 62
rect -321 -100 -255 -62
rect -225 62 -159 100
rect -225 -62 -209 62
rect -175 -62 -159 62
rect -225 -100 -159 -62
rect -129 62 -63 100
rect -129 -62 -113 62
rect -79 -62 -63 62
rect -129 -100 -63 -62
rect -33 62 33 100
rect -33 -62 -17 62
rect 17 -62 33 62
rect -33 -100 33 -62
rect 63 62 129 100
rect 63 -62 79 62
rect 113 -62 129 62
rect 63 -100 129 -62
rect 159 62 225 100
rect 159 -62 175 62
rect 209 -62 225 62
rect 159 -100 225 -62
rect 255 62 321 100
rect 255 -62 271 62
rect 305 -62 321 62
rect 255 -100 321 -62
rect 351 74 409 100
rect 351 62 413 74
rect 351 -62 367 62
rect 401 -62 413 62
rect 351 -74 413 -62
rect 351 -100 409 -74
<< ndiffc >>
rect -401 -62 -367 62
rect -305 -62 -271 62
rect -209 -62 -175 62
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
rect 175 -62 209 62
rect 271 -62 305 62
rect 367 -62 401 62
<< poly >>
rect -351 100 -321 136
rect -255 100 -225 136
rect -159 100 -129 134
rect -63 100 -33 134
rect 33 100 63 134
rect 129 100 159 134
rect 225 100 255 136
rect 321 100 351 134
rect -351 -120 -321 -100
rect -255 -120 -225 -100
rect -159 -120 -129 -100
rect -63 -120 -33 -100
rect 33 -120 63 -100
rect 129 -120 159 -100
rect 225 -120 255 -100
rect 321 -120 351 -100
rect -353 -162 351 -120
<< locali >>
rect 321 116 351 134
rect -401 62 -367 78
rect -401 -78 -367 -62
rect -305 62 -271 78
rect -305 -78 -271 -62
rect -209 62 -175 78
rect -209 -78 -175 -62
rect -113 62 -79 78
rect -113 -78 -79 -62
rect -17 62 17 78
rect -17 -78 17 -62
rect 79 62 113 78
rect 79 -78 113 -62
rect 175 62 209 78
rect 175 -78 209 -62
rect 271 62 305 78
rect 271 -78 305 -62
rect 367 62 401 78
rect 367 -78 401 -62
<< viali >>
rect -401 -62 -367 62
rect -305 -62 -271 62
rect -209 -62 -175 62
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
rect 175 -62 209 62
rect 271 -62 305 62
rect 367 -62 401 62
<< metal1 >>
rect -407 62 -361 74
rect -407 -62 -401 62
rect -367 -62 -361 62
rect -407 -74 -361 -62
rect -311 62 -265 74
rect -311 -62 -305 62
rect -271 -62 -265 62
rect -311 -74 -265 -62
rect -215 62 -169 74
rect -215 -62 -209 62
rect -175 -62 -169 62
rect -215 -74 -169 -62
rect -119 62 -73 74
rect -119 -62 -113 62
rect -79 -62 -73 62
rect -119 -74 -73 -62
rect -23 62 23 74
rect -23 -62 -17 62
rect 17 -62 23 62
rect -23 -74 23 -62
rect 73 62 119 74
rect 73 -62 79 62
rect 113 -62 119 62
rect 73 -74 119 -62
rect 169 62 215 74
rect 169 -62 175 62
rect 209 -62 215 62
rect 169 -74 215 -62
rect 265 62 311 74
rect 265 -62 271 62
rect 305 -62 311 62
rect 265 -74 311 -62
rect 361 62 407 74
rect 361 -62 367 62
rect 401 -62 407 62
rect 361 -74 407 -62
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.150 m 1 nf 8 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
