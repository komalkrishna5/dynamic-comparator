magic
tech sky130A
magscale 1 2
timestamp 1646324451
<< error_p >>
rect -261 174 -227 224
rect -209 140 -203 192
rect 195 140 209 192
rect 229 174 263 224
rect -261 -290 -225 -234
rect -261 -726 -223 -674
rect 225 -726 263 -674
<< nwell >>
rect -261 -210 263 200
<< pmos >>
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
<< pdiff >>
rect -217 74 -159 100
rect -221 62 -159 74
rect -221 -62 -209 62
rect -175 -62 -159 62
rect -221 -74 -159 -62
rect -217 -100 -159 -74
rect -129 62 -63 100
rect -129 -62 -113 62
rect -79 -62 -63 62
rect -129 -100 -63 -62
rect -33 62 33 100
rect -33 -62 -17 62
rect 17 -62 33 62
rect -33 -100 33 -62
rect 63 62 129 100
rect 63 -62 79 62
rect 113 -62 129 62
rect 63 -100 129 -62
rect 159 74 217 100
rect 159 62 221 74
rect 159 -62 175 62
rect 209 -62 221 62
rect 159 -74 221 -62
rect 159 -100 217 -74
<< pdiffc >>
rect -209 -62 -175 62
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
rect 175 -62 209 62
<< poly >>
rect -159 100 -129 138
rect -63 100 -33 138
rect 33 100 63 138
rect 129 100 159 138
rect -159 -120 -129 -100
rect -63 -120 -33 -100
rect 33 -120 63 -100
rect 129 -120 159 -100
rect -159 -152 161 -120
rect 15 -208 45 -152
<< locali >>
rect -261 174 -237 224
rect -209 62 -175 192
rect -209 -78 -175 -62
rect -113 62 -79 78
rect -113 -68 -79 -62
rect -115 -116 -79 -68
rect -17 62 17 192
rect -17 -78 17 -62
rect 79 62 113 78
rect 79 -64 113 -62
rect 77 -116 113 -64
rect 175 62 209 192
rect 229 174 263 224
rect 175 -78 209 -62
rect -115 -154 113 -116
rect 61 -220 95 -154
rect -261 -290 -225 -234
rect 217 -290 263 -234
rect -261 -726 -223 -674
rect 225 -726 263 -674
<< viali >>
rect -209 -62 -175 62
rect -113 -62 -79 62
rect -17 -62 17 62
rect 79 -62 113 62
rect 175 -62 209 62
<< metal1 >>
rect -215 62 -169 74
rect -215 -62 -209 62
rect -175 -62 -169 62
rect -215 -74 -169 -62
rect -119 62 -73 74
rect -119 -62 -113 62
rect -79 -62 -73 62
rect -119 -74 -73 -62
rect -23 62 23 74
rect -23 -62 -17 62
rect 17 -62 23 62
rect -23 -74 23 -62
rect 73 62 119 74
rect 73 -62 79 62
rect 113 -62 119 62
rect 73 -74 119 -62
rect 169 62 215 74
rect 169 -62 175 62
rect 209 -62 215 62
rect 169 -74 215 -62
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 4 diffcov 70 polycov 70 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 70 rlcov 70 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 70 viadrn 70 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
