magic
tech sky130A
timestamp 1646599058
<< poly >>
rect 263 2110 303 2122
rect 263 2093 273 2110
rect 290 2107 303 2110
rect 364 2107 379 2121
rect 661 2110 701 2122
rect 661 2108 671 2110
rect 290 2093 379 2107
rect 263 2091 379 2093
rect 562 2093 671 2108
rect 688 2093 701 2110
rect 562 2092 701 2093
rect 263 2080 303 2091
rect 661 2080 701 2092
<< polycont >>
rect 273 2093 290 2110
rect 671 2093 688 2110
<< locali >>
rect 263 2110 298 2118
rect 263 2093 273 2110
rect 290 2093 298 2110
rect 263 2089 298 2093
rect 661 2110 696 2118
rect 661 2093 671 2110
rect 688 2093 696 2110
rect 661 2089 696 2093
rect 823 1514 851 1564
rect 823 1497 828 1514
rect 846 1497 851 1514
rect 823 1496 851 1497
<< viali >>
rect 153 1539 178 1562
rect 692 1539 717 1562
rect 828 1497 846 1514
<< metal1 >>
rect 263 2113 303 2122
rect -104 2087 303 2113
rect -104 1564 -64 2087
rect 263 2080 303 2087
rect 661 2116 701 2122
rect 661 2089 986 2116
rect 661 2080 701 2089
rect 136 1564 187 1572
rect -104 1562 187 1564
rect -104 1539 153 1562
rect 178 1539 187 1562
rect -104 1536 187 1539
rect -104 199 -64 1536
rect 136 1515 187 1536
rect 684 1562 726 1572
rect 684 1539 692 1562
rect 717 1561 726 1562
rect 946 1561 986 2089
rect 717 1539 987 1561
rect 684 1536 987 1539
rect 684 1530 726 1536
rect 823 1515 852 1520
rect 136 1514 852 1515
rect 136 1497 828 1514
rect 846 1497 852 1514
rect 946 1501 987 1536
rect 136 1496 852 1497
rect 823 1490 852 1496
rect -29 965 153 996
rect 601 969 903 1000
rect -29 293 -1 965
rect 130 950 153 965
rect 130 944 152 950
rect 875 293 903 969
rect -29 272 20 293
rect 858 272 903 293
rect 947 206 987 1501
rect -104 171 35 199
rect 819 178 987 206
use SR_latch  SR_latch_0 ~/mycomparator_copy1/layout/latch
timestamp 1646507701
transform 1 0 235 0 1 2046
box 0 0 436 474
use latch_2  latch_2_0 ~/mycomparator_copy1/layout/latch
timestamp 1646503715
transform 1 0 43 0 1 1318
box 0 0 801 501
use preamp_part1  preamp_part1_0 ~/mycomparator_copy1/layout/preamp
timestamp 1646568821
transform 1 0 360 0 1 130
box -360 -130 510 508
use preamp_part2  preamp_part2_0 ~/mycomparator_copy1/layout/preamp
timestamp 1646595273
transform 1 0 69 0 1 688
box 58 1 641 544
<< end >>
