* SPICE3 file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_AC5Z8B a_159_n100# li_217_n290# li_n261_n290# li_229_174#
+ a_n221_n74# a_n129_n100# a_n159_n152# li_225_n726# a_n33_n100# w_n261_n210# li_n261_174#
+ li_n261_n726# VSUBS
X0 a_n129_n100# a_n159_n152# a_n33_n100# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=5.32e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n159_n152# a_n129_n100# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_159_n100# a_n159_n152# a_n129_n100# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_n129_n100# a_n159_n152# a_n221_n74# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_XJTKXQ a_33_n122# a_n63_n122# a_63_n100# a_n125_n74#
+ a_n33_n100# VSUBS
X0 a_63_n100# a_33_n122# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n122# a_n125_n74# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt inv_W2 sky130_fd_pr__pfet_01v8_AC5Z8B_0/w_n261_n210# Vout Vin VDD GND VSUBS
Xsky130_fd_pr__pfet_01v8_AC5Z8B_0 VDD Vout Vin VDD VDD Vout Vin GND VDD sky130_fd_pr__pfet_01v8_AC5Z8B_0/w_n261_n210#
+ VDD GND VSUBS sky130_fd_pr__pfet_01v8_AC5Z8B
Xsky130_fd_pr__nfet_01v8_XJTKXQ_0 Vin Vin GND GND Vout VSUBS sky130_fd_pr__nfet_01v8_XJTKXQ
.ends

.subckt sky130_fd_pr__nfet_01v8_7RYEVP a_n73_n69# a_n33_n157# a_15_n69# VSUBS
X0 a_15_n69# a_n33_n157# a_n73_n69# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt nmos_1u sky130_fd_pr__nfet_01v8_7RYEVP_0/VSUBS sky130_fd_pr__nfet_01v8_7RYEVP_0/a_15_n69#
+ m1_n86_2#
Xsky130_fd_pr__nfet_01v8_7RYEVP_0 sky130_fd_pr__nfet_01v8_7RYEVP_0/VSUBS m1_n86_2#
+ sky130_fd_pr__nfet_01v8_7RYEVP_0/a_15_n69# sky130_fd_pr__nfet_01v8_7RYEVP_0/VSUBS
+ sky130_fd_pr__nfet_01v8_7RYEVP
.ends

.subckt pmos_2uf2 a_63_n100# a_33_n130# w_n317_n202# a_n33_n100# a_n63_n130# VSUBS
X0 a_63_n100# a_33_n130# a_n33_n100# w_n317_n202# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n130# w_n317_n202# w_n317_n202# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.8e+11p ps=2.76e+06u w=1e+06u l=150000u
.ends

.subckt inv_W1 Vout VDD Vin GND
Xnmos_1u_0 GND Vout Vin nmos_1u
Xpmos_2uf2_0 VDD Vin VDD Vout Vin GND pmos_2uf2
.ends

.subckt buffer_1#0 inv_W2_0/VDD inv_W2_0/Vout inv_W1_0/Vin VSUBS
Xinv_W2_0 inv_W2_0/VDD inv_W2_0/Vout inv_W2_0/Vin inv_W2_0/VDD VSUBS VSUBS inv_W2
Xinv_W1_0 inv_W2_0/Vin inv_W2_0/VDD inv_W1_0/Vin VSUBS inv_W1
.ends

.subckt buffer_1 inv_W2_0/VDD inv_W2_0/Vout inv_W1_0/Vin inv_W2_0/Vin VSUBS
Xinv_W2_0 inv_W2_0/VDD inv_W2_0/Vout inv_W2_0/Vin inv_W2_0/VDD VSUBS VSUBS inv_W2
Xinv_W1_0 inv_W2_0/Vin inv_W2_0/VDD inv_W1_0/Vin VSUBS inv_W1
.ends

.subckt sky130_fd_pr__nfet_01v8_KZU588 a_159_n100# a_255_n100# a_351_n100# a_n129_n100#
+ a_63_n100# li_321_116# a_n353_n162# a_n225_n100# a_n413_n74# a_n321_n100# a_n33_n100#
+ VSUBS
X0 a_n321_n100# a_n353_n162# a_n413_n74# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
X1 a_n225_n100# a_n353_n162# a_n321_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_n129_n100# a_n353_n162# a_n225_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_63_n100# a_n353_n162# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 a_n33_n100# a_n353_n162# a_n129_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_351_n100# a_n353_n162# a_255_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6 a_159_n100# a_n353_n162# a_63_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_255_n100# a_n353_n162# a_159_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_RL4NCG a_543_n100# a_159_n100# a_n609_n100# a_321_n126#
+ a_n705_n100# a_255_n100# a_n159_n128# a_n543_n128# a_n255_n126# a_351_n100# a_n417_n100#
+ a_33_n128# a_n129_n100# a_n513_n100# a_n351_n128# a_63_n100# w_n833_n200# a_n225_n100#
+ a_609_n128# a_n63_n126# a_n797_n74# a_705_n126# a_n321_n100# a_639_n100# a_417_n128#
+ a_n639_n126# a_735_n100# a_n33_n100# a_513_n126# a_129_n126# a_447_n100# a_n735_n128#
+ a_n447_n126# a_225_n128# VSUBS
X0 a_63_n100# a_33_n128# a_n33_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n126# a_n129_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_255_n100# a_225_n128# a_159_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_351_n100# a_321_n126# a_255_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_543_n100# a_513_n126# a_447_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X5 a_159_n100# a_129_n126# a_63_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_447_n100# a_417_n128# a_351_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_639_n100# a_609_n128# a_543_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_735_n100# a_705_n126# a_639_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_n513_n100# a_n543_n128# a_n609_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10 a_n321_n100# a_n351_n128# a_n417_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X11 a_n225_n100# a_n255_n126# a_n321_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_n705_n100# a_n735_n128# a_n797_n74# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
X13 a_n609_n100# a_n639_n126# a_n705_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_n417_n100# a_n447_n126# a_n513_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_n129_n100# a_n159_n128# a_n225_n100# w_n833_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt inv_W8 li_354_902# w_354_500# li_354_0# li_512_546# a_804_430# VSUBS
Xsky130_fd_pr__nfet_01v8_KZU588_0 li_354_0# li_512_546# li_354_0# li_512_546# li_512_546#
+ li_512_546# a_804_430# li_354_0# li_354_0# li_512_546# li_354_0# VSUBS sky130_fd_pr__nfet_01v8_KZU588
Xsky130_fd_pr__pfet_01v8_RL4NCG_0 li_354_902# li_354_902# li_354_902# a_804_430# li_512_546#
+ li_512_546# a_804_430# a_804_430# a_804_430# li_354_902# li_354_902# a_804_430#
+ li_512_546# li_512_546# a_804_430# li_512_546# w_354_500# li_354_902# a_804_430#
+ a_804_430# li_354_902# a_804_430# li_512_546# li_512_546# a_804_430# a_804_430#
+ li_354_902# li_354_902# a_804_430# a_804_430# li_512_546# a_804_430# a_804_430#
+ a_804_430# VSUBS sky130_fd_pr__pfet_01v8_RL4NCG
.ends

.subckt sky130_fd_pr__nfet_01v8_VJWT33 a_543_n100# a_159_n100# a_n609_n100# a_n705_n100#
+ a_255_n100# a_351_n100# a_n417_n100# a_n129_n100# a_n513_n100# a_63_n100# a_n225_n100#
+ a_n797_n74# a_n735_n176# a_n321_n100# a_639_n100# a_735_n100# a_n33_n100# a_447_n100#
+ VSUBS
X0 a_n513_n100# a_n735_n176# a_n609_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n321_n100# a_n735_n176# a_n417_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_n225_n100# a_n735_n176# a_n321_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_n705_n100# a_n735_n176# a_n797_n74# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
X4 a_n609_n100# a_n735_n176# a_n705_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_n417_n100# a_n735_n176# a_n513_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_n129_n100# a_n735_n176# a_n225_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_63_n100# a_n735_n176# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X8 a_n33_n100# a_n735_n176# a_n129_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_351_n100# a_n735_n176# a_255_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10 a_159_n100# a_n735_n176# a_63_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_255_n100# a_n735_n176# a_159_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_447_n100# a_n735_n176# a_351_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X13 a_543_n100# a_n735_n176# a_447_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_639_n100# a_n735_n176# a_543_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_735_n100# a_n735_n176# a_639_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_3M44SC a_543_n100# a_159_n100# a_n609_n100# a_321_n126#
+ a_1473_n126# a_1089_n126# a_n1407_n126# a_n705_n100# a_255_n100# a_n159_n128# a_n543_n128#
+ a_1407_n100# a_1185_n128# a_n255_n126# a_351_n100# a_n417_n100# a_n801_n100# a_n1119_n128#
+ a_n1503_n128# a_1281_n126# a_897_n126# a_33_n128# w_n1601_n200# a_1503_n100# a_1119_n100#
+ a_n1377_n100# a_n1215_n126# a_n129_n100# a_n513_n100# a_n351_n128# a_n1565_n74#
+ a_1215_n100# a_63_n100# a_n1089_n100# a_n1473_n100# a_993_n128# a_n225_n100# a_609_n128#
+ a_n63_n126# a_n1311_n128# a_1311_n100# a_927_n100# a_n1185_n100# a_705_n126# a_n1023_n126#
+ a_n321_n100# a_1023_n100# a_639_n100# a_n1281_n100# a_n927_n128# a_801_n128# a_417_n128#
+ a_n639_n126# a_735_n100# a_n33_n100# a_513_n126# a_129_n126# a_n897_n100# a_831_n100#
+ a_447_n100# a_n735_n128# a_n993_n100# a_n447_n126# a_n831_n126# a_1377_n128# a_225_n128#
+ VSUBS
X0 a_63_n100# a_33_n128# a_n33_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_927_n100# a_897_n126# a_831_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_1023_n100# a_993_n128# a_927_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_1311_n100# a_1281_n126# a_1215_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 a_1119_n100# a_1089_n126# a_1023_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_1215_n100# a_1185_n128# a_1119_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_1407_n100# a_1377_n128# a_1311_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_1503_n100# a_1473_n126# a_1407_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_n33_n100# a_n63_n126# a_n129_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X9 a_255_n100# a_225_n128# a_159_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10 a_351_n100# a_321_n126# a_255_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_543_n100# a_513_n126# a_447_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X12 a_831_n100# a_801_n128# a_735_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X13 a_159_n100# a_129_n126# a_63_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_447_n100# a_417_n128# a_351_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_639_n100# a_609_n128# a_543_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X16 a_735_n100# a_705_n126# a_639_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_n1281_n100# a_n1311_n128# a_n1377_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X18 a_n993_n100# a_n1023_n126# a_n1089_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X19 a_n1473_n100# a_n1503_n128# a_n1565_n74# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
X20 a_n1377_n100# a_n1407_n126# a_n1473_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_n1185_n100# a_n1215_n126# a_n1281_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X22 a_n1089_n100# a_n1119_n128# a_n1185_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_n801_n100# a_n831_n126# a_n897_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X24 a_n513_n100# a_n543_n128# a_n609_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X25 a_n321_n100# a_n351_n128# a_n417_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X26 a_n225_n100# a_n255_n126# a_n321_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X27 a_n897_n100# a_n927_n128# a_n993_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n705_n100# a_n735_n128# a_n801_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X29 a_n609_n100# a_n639_n126# a_n705_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_n417_n100# a_n447_n126# a_n513_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_n129_n100# a_n159_n128# a_n225_n100# w_n1601_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
C0 w_n1601_n200# VSUBS 3.82fF
.ends

.subckt inv_W16 li_128_546# li_n14_902# a_82_816# w_82_814# li_n14_0# VSUBS
Xsky130_fd_pr__nfet_01v8_VJWT33_0 li_n14_0# li_n14_0# li_n14_0# li_128_546# li_128_546#
+ li_n14_0# li_n14_0# li_128_546# li_128_546# li_128_546# li_n14_0# li_n14_0# a_82_816#
+ li_128_546# li_128_546# li_n14_0# li_n14_0# li_128_546# VSUBS sky130_fd_pr__nfet_01v8_VJWT33
Xsky130_fd_pr__pfet_01v8_3M44SC_0 li_n14_902# li_n14_902# li_n14_902# a_82_816# a_82_816#
+ a_82_816# a_82_816# li_128_546# li_128_546# a_82_816# a_82_816# li_128_546# a_82_816#
+ a_82_816# li_n14_902# li_n14_902# li_n14_902# a_82_816# a_82_816# a_82_816# a_82_816#
+ a_82_816# w_82_814# li_n14_902# li_n14_902# li_n14_902# a_82_816# li_128_546# li_128_546#
+ a_82_816# li_n14_902# li_128_546# li_128_546# li_128_546# li_128_546# a_82_816#
+ li_n14_902# a_82_816# a_82_816# a_82_816# li_n14_902# li_n14_902# li_n14_902# a_82_816#
+ a_82_816# li_128_546# li_128_546# li_128_546# li_128_546# a_82_816# a_82_816# a_82_816#
+ a_82_816# li_n14_902# li_n14_902# a_82_816# a_82_816# li_128_546# li_128_546# li_128_546#
+ a_82_816# li_n14_902# a_82_816# a_82_816# a_82_816# a_82_816# VSUBS sky130_fd_pr__pfet_01v8_3M44SC
C0 a_82_816# VSUBS 2.90fF
C1 w_82_814# VSUBS 3.92fF
.ends

.subckt buffer_2 Vout inv_W8_0/li_354_902# w_1666_500# inv_W8_0/a_804_430# inv_W8_0/li_354_0#
+ VSUBS
Xinv_W8_0 inv_W8_0/li_354_902# w_1666_500# inv_W8_0/li_354_0# inv_W16_0/a_82_816#
+ inv_W8_0/a_804_430# VSUBS inv_W8
Xinv_W16_0 Vout inv_W8_0/li_354_902# inv_W16_0/a_82_816# w_1666_500# inv_W8_0/li_354_0#
+ VSUBS inv_W16
C0 inv_W8_0/li_354_902# VSUBS -3.18fF
C1 w_1666_500# VSUBS 6.52fF
C2 inv_W8_0/li_354_0# VSUBS 2.10fF
.ends

.subckt buffer_12 buffer_1_0/inv_W2_0/Vout buf_in buffer_1_0/inv_W2_0/Vin VDD buf_out
+ GND
Xbuffer_1_0 VDD buffer_1_0/inv_W2_0/Vout buf_in buffer_1_0/inv_W2_0/Vin GND buffer_1
Xbuffer_2_0 buf_out VDD VDD buffer_1_0/inv_W2_0/Vout GND GND buffer_2
C0 VDD 0 3.98fF
C1 GND 0 2.58fF
.ends

.subckt sky130_fd_pr__pfet_01v8_RFM3CD a_n73_n100# w_n109_n162# a_15_n100# a_n15_n126#
+ VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# w_n109_n162# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_F5U58G#0 a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_XJTKXQ#0 a_n63_n152# a_63_n100# a_n125_n74# a_n33_n100#
+ VSUBS
X0 a_63_n100# a_n63_n152# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n152# a_n125_n74# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt preamp_part2 a_148_644# sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126# a_380_480#
+ sky130_fd_pr__pfet_01v8_RFM3CD_1/w_n109_n162# sky130_fd_pr__pfet_01v8_RFM3CD_0/a_n15_n126#
+ sky130_fd_pr__pfet_01v8_RFM3CD_1/a_n15_n126# a_1170_652# sky130_fd_pr__pfet_01v8_RFM3CD_0/w_n109_n162#
+ VDD GND a_792_2# VSUBS
Xsky130_fd_pr__pfet_01v8_RFM3CD_0 VDD sky130_fd_pr__pfet_01v8_RFM3CD_0/w_n109_n162#
+ li_210_488# sky130_fd_pr__pfet_01v8_RFM3CD_0/a_n15_n126# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD
Xsky130_fd_pr__pfet_01v8_RFM3CD_1 li_928_394# sky130_fd_pr__pfet_01v8_RFM3CD_1/w_n109_n162#
+ VDD sky130_fd_pr__pfet_01v8_RFM3CD_1/a_n15_n126# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD
Xsky130_fd_pr__nfet_01v8_F5U58G_0 m1_322_206# GND sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126#
+ VSUBS sky130_fd_pr__nfet_01v8_F5U58G#0
Xsky130_fd_pr__nfet_01v8_F5U58G_1 a_792_2# li_210_488# a_148_644# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#0
Xsky130_fd_pr__nfet_01v8_F5U58G_2 li_928_394# a_380_480# a_1170_652# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#0
Xsky130_fd_pr__nfet_01v8_XJTKXQ_0 a_380_480# m1_322_206# m1_322_206# li_210_488# VSUBS
+ sky130_fd_pr__nfet_01v8_XJTKXQ#0
Xsky130_fd_pr__nfet_01v8_XJTKXQ_1 a_792_2# m1_322_206# m1_322_206# li_928_394# VSUBS
+ sky130_fd_pr__nfet_01v8_XJTKXQ#0
.ends

.subckt sky130_fd_pr__nfet_01v8_F5U58G a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_AC5E9B w_n161_n200# a_33_n126# a_63_n100# a_n125_n74#
+ a_n33_n100# a_n63_n130# VSUBS
X0 a_63_n100# a_33_n126# a_n33_n100# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n130# a_n125_n74# w_n161_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt SR_latch a_648_848# sky130_fd_pr__nfet_01v8_F5U58G_1/a_n15_n126# sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126#
+ a_262_508# VDD w_0_524# GND VSUBS
Xsky130_fd_pr__nfet_01v8_F5U58G_0 a_648_848# GND sky130_fd_pr__nfet_01v8_F5U58G_0/a_n15_n126#
+ VSUBS sky130_fd_pr__nfet_01v8_F5U58G
Xsky130_fd_pr__nfet_01v8_F5U58G_1 GND a_262_508# sky130_fd_pr__nfet_01v8_F5U58G_1/a_n15_n126#
+ VSUBS sky130_fd_pr__nfet_01v8_F5U58G
Xsky130_fd_pr__pfet_01v8_AC5E9B_0 w_0_524# a_262_508# VDD VDD a_648_848# a_262_508#
+ VSUBS sky130_fd_pr__pfet_01v8_AC5E9B
Xsky130_fd_pr__pfet_01v8_AC5E9B_1 w_0_524# a_648_848# VDD VDD a_262_508# a_648_848#
+ VSUBS sky130_fd_pr__pfet_01v8_AC5E9B
.ends

.subckt sky130_fd_pr__nfet_01v8_G6PLX8 a_159_n100# a_n221_n74# a_n129_n100# a_63_n100#
+ a_n33_n100# a_n159_n122# VSUBS
X0 a_n129_n100# a_n159_n122# a_n221_n74# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
X1 a_63_n100# a_n159_n122# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_n33_n100# a_n159_n122# a_n129_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_159_n100# a_n159_n122# a_63_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_F5U58G#1 a_n73_n100# a_15_n100# a_n15_n126# VSUBS
X0 a_15_n100# a_n15_n126# a_n73_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_8FHE5N a_n33_n50# a_63_n50# a_n63_n76# a_33_n76# a_n125_n39#
+ VSUBS
X0 a_n33_n50# a_n63_n76# a_n125_n39# VSUBS sky130_fd_pr__nfet_01v8 ad=1.65e+11p pd=1.66e+06u as=1.528e+11p ps=1.62e+06u w=500000u l=150000u
X1 a_63_n50# a_33_n76# a_n33_n50# VSUBS sky130_fd_pr__nfet_01v8 ad=1.528e+11p pd=1.62e+06u as=0p ps=0u w=500000u l=150000u
.ends

.subckt preamp_part1 li_954_42# li_n718_44# a_n656_268# a_80_n258# a_n302_940# w_n720_482#
+ a_n434_n260# a_506_940# a_864_270# VDD a_388_n260# GND VSUBS
Xsky130_fd_pr__nfet_01v8_G6PLX8_0 li_n484_188# li_n484_188# a_n656_268# a_n656_268#
+ li_n484_188# a_n434_n260# VSUBS sky130_fd_pr__nfet_01v8_G6PLX8
Xsky130_fd_pr__nfet_01v8_G6PLX8_1 li_n484_188# li_n484_188# a_864_270# a_864_270#
+ li_n484_188# a_388_n260# VSUBS sky130_fd_pr__nfet_01v8_G6PLX8
Xsky130_fd_pr__pfet_01v8_RFM3CD_0 VDD w_n720_482# a_n656_268# a_n302_940# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD
Xsky130_fd_pr__pfet_01v8_RFM3CD_1 a_864_270# w_n720_482# VDD a_506_940# VSUBS sky130_fd_pr__pfet_01v8_RFM3CD
Xsky130_fd_pr__nfet_01v8_F5U58G_0 li_n718_44# GND a_n656_268# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#1
Xsky130_fd_pr__nfet_01v8_F5U58G_1 GND li_954_42# a_864_270# VSUBS sky130_fd_pr__nfet_01v8_F5U58G#1
Xsky130_fd_pr__nfet_01v8_8FHE5N_0 li_n484_188# GND a_80_n258# a_80_n258# GND VSUBS
+ sky130_fd_pr__nfet_01v8_8FHE5N
.ends

.subckt sky130_fd_pr__pfet_01v8_AC5Z8B#0 a_159_n100# li_217_n290# li_n261_n290# li_229_174#
+ a_n221_n74# a_n129_n100# a_n159_n152# li_225_n726# a_n33_n100# w_n261_n210# li_n261_174#
+ li_n261_n726# VSUBS
X0 a_n129_n100# a_n159_n152# a_n33_n100# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=6.6e+11p pd=5.32e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n159_n152# a_n129_n100# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_159_n100# a_n159_n152# a_n129_n100# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=3.048e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_n129_n100# a_n159_n152# a_n221_n74# w_n261_n210# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_XJTKXQ#1 a_33_n122# a_n63_n122# a_63_n100# a_n125_n74#
+ a_n33_n100# VSUBS
X0 a_63_n100# a_33_n122# a_n33_n100# VSUBS sky130_fd_pr__nfet_01v8 ad=3.048e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n63_n122# a_n125_n74# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.048e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt inv_W2#0 sky130_fd_pr__pfet_01v8_AC5Z8B_0/w_n261_n210# Vout Vin VDD GND VSUBS
Xsky130_fd_pr__pfet_01v8_AC5Z8B_0 VDD Vout Vin VDD VDD Vout Vin GND VDD sky130_fd_pr__pfet_01v8_AC5Z8B_0/w_n261_n210#
+ VDD GND VSUBS sky130_fd_pr__pfet_01v8_AC5Z8B#0
Xsky130_fd_pr__nfet_01v8_XJTKXQ_0 Vin Vin GND GND Vout VSUBS sky130_fd_pr__nfet_01v8_XJTKXQ#1
.ends

.subckt sky130_fd_pr__pfet_01v8_5SVZDE a_n111_n158# a_n173_n100# a_15_n100# a_111_n100#
+ a_n81_n100# w_n789_n196# VSUBS
X0 a_15_n100# a_n111_n158# a_n81_n100# w_n789_n196# sky130_fd_pr__pfet_01v8 ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_111_n100# a_n111_n158# a_15_n100# w_n789_n196# sky130_fd_pr__pfet_01v8 ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_n81_n100# a_n111_n158# a_n173_n100# w_n789_n196# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt latch_2 m1_718_782# inv_W2_1/Vin inv_W2_1/GND sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196#
+ sky130_fd_pr__pfet_01v8_5SVZDE_0/a_n111_n158# inv_W2_0/Vin inv_W2_1/Vout VSUBS
Xinv_W2_0 sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196# inv_W2_1/Vin inv_W2_0/Vin
+ inv_W2_1/VDD inv_W2_1/GND VSUBS inv_W2#0
Xinv_W2_1 sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196# inv_W2_1/Vout inv_W2_1/Vin
+ inv_W2_1/VDD inv_W2_1/GND VSUBS inv_W2#0
Xsky130_fd_pr__pfet_01v8_5SVZDE_0 sky130_fd_pr__pfet_01v8_5SVZDE_0/a_n111_n158# inv_W2_1/VDD
+ inv_W2_1/VDD m1_718_782# m1_718_782# sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196#
+ VSUBS sky130_fd_pr__pfet_01v8_5SVZDE
C0 sky130_fd_pr__pfet_01v8_5SVZDE_0/w_n789_n196# VSUBS 2.01fF
.ends

.subckt compaartor_v4 Outn Vp Vn CLK VDD GND Outp CLKBAR
Xpreamp_part2_0 CLK CLK m1_1202_1938# VDD CLK CLK CLK VDD VDD GND m1_n58_544# GND
+ preamp_part2
XSR_latch_0 Outp latch_2_0/inv_W2_1/Vin latch_2_0/inv_W2_0/Vin Outn VDD VDD GND GND
+ SR_latch
Xpreamp_part1_0 latch_2_0/inv_W2_1/Vin latch_2_0/inv_W2_0/Vin m1_n58_544# CLK CLK
+ VDD Vn CLK m1_1202_1938# VDD Vp GND GND preamp_part1
Xlatch_2_0 VDD latch_2_0/inv_W2_1/Vin GND VDD CLKBAR latch_2_0/inv_W2_0/Vin latch_2_0/inv_W2_0/Vin
+ GND latch_2
C0 latch_2_0/inv_W2_1/Vin GND 2.84fF
C1 latch_2_0/inv_W2_0/Vin GND 4.28fF
C2 CLK GND 17.54fF
C3 VDD GND 22.81fF
C4 m1_n58_544# GND 2.08fF
.ends

.subckt buffer_2#0 Vout w_1666_500# inv_W8_0/li_354_902# inv_W8_0/a_804_430# inv_W8_0/li_354_0#
+ VSUBS
Xinv_W8_0 inv_W8_0/li_354_902# w_1666_500# inv_W8_0/li_354_0# inv_W16_0/a_82_816#
+ inv_W8_0/a_804_430# VSUBS inv_W8
Xinv_W16_0 Vout inv_W8_0/li_354_902# inv_W16_0/a_82_816# w_1666_500# inv_W8_0/li_354_0#
+ VSUBS inv_W16
C0 inv_W8_0/li_354_902# VSUBS -3.18fF
C1 w_1666_500# VSUBS 6.52fF
C2 inv_W8_0/li_354_0# VSUBS 2.10fF
.ends

.subckt buffer_2#1 Vout w_1666_500# inv_W8_0/li_354_902# inv_W8_0/a_804_430# inv_W8_0/li_354_0#
+ VSUBS
Xinv_W8_0 inv_W8_0/li_354_902# w_1666_500# inv_W8_0/li_354_0# inv_W16_0/a_82_816#
+ inv_W8_0/a_804_430# VSUBS inv_W8
Xinv_W16_0 Vout inv_W8_0/li_354_902# inv_W16_0/a_82_816# w_1666_500# inv_W8_0/li_354_0#
+ VSUBS inv_W16
C0 inv_W8_0/li_354_902# VSUBS -3.18fF
C1 w_1666_500# VSUBS 6.52fF
C2 inv_W8_0/li_354_0# VSUBS 2.10fF
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[5] io_analog[6] io_analog[7] io_analog[8]
+ io_analog[9] io_analog[4] io_clamp_high[0] io_clamp_low[0] io_in[0] io_in[10] io_in[11]
+ io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19]
+ io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10]
+ io_in_3v3[11] io_in_3v3[12] io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16]
+ io_in_3v3[17] io_in_3v3[18] io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21]
+ io_in_3v3[22] io_in_3v3[23] io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2]
+ io_in_3v3[3] io_in_3v3[4] io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9]
+ io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16]
+ io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23]
+ io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6]
+ io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13]
+ io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20]
+ io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xbuffer_1_0 vccd1 L1 compaartor_v4_0/Outn vssa1 buffer_1#0
Xbuffer_1_1 vccd1 L2 compaartor_v4_0/Outp vssa1 buffer_1#0
Xbuffer_12_0 L4 io_analog[8] L3 vccd1 compaartor_v4_0/CLK vssa1 buffer_12
Xbuffer_12_1 buffer_12_1/buffer_1_0/inv_W2_0/Vout io_analog[7] buffer_12_1/buffer_1_0/inv_W2_0/Vin
+ vccd1 CB vssa1 buffer_12
Xcompaartor_v4_0 compaartor_v4_0/Outn io_analog[5] io_analog[6] compaartor_v4_0/CLK
+ vccd1 vssa1 compaartor_v4_0/Outp CB compaartor_v4
Xbuffer_2_0 io_analog[3] vccd1 vccd1 L1 vssa1 vssa1 buffer_2#0
Xbuffer_2_1 io_analog[2] vccd1 vccd1 L2 vssa1 vssa1 buffer_2#1
C0 m4_204098_586508# io_analog[5] 518.20fF
C1 vccd1 m4_186716_584374# 104.50fF
C2 CB io_analog[5] 3.06fF
C3 vccd1 io_analog[2] 35.31fF
C4 vccd1 io_analog[5] 42.19fF
C5 vccd1 io_analog[6] 40.88fF
C6 io_analog[7] m4_186716_584374# 4.20fF
C7 vccd1 m4_204098_586508# 119.00fF
C8 vccd1 compaartor_v4_0/Outn 67.00fF
C9 io_analog[5] io_analog[7] 75.42fF
C10 m4_204098_586508# io_analog[7] 4.77fF
C11 m4_186716_584374# io_analog[8] 4.20fF
C12 io_analog[6] compaartor_v4_0/CLK 2.02fF
C13 io_analog[3] vccd1 35.18fF
C14 m3_417434_589490# vccd1 7.13fF
C15 CB compaartor_v4_0/CLK 3.22fF
C16 io_analog[6] m4_186716_584374# 469.66fF
C17 vccd1 compaartor_v4_0/Outp 66.83fF
C18 io_analog[4] vssa1 25.05fF
C19 vssd2 vssa1 13.04fF
C20 vssd1 vssa1 13.62fF
C21 vdda2 vssa1 13.04fF
C22 vdda1 vssa1 26.08fF
C23 vssa2 vssa1 13.04fF
C24 io_analog[0] vssa1 6.83fF
C25 io_analog[1] vssa1 6.83fF
C26 io_clamp_high[0] vssa1 3.58fF
C27 io_clamp_low[0] vssa1 3.58fF
C28 vccd2 vssa1 13.04fF
C29 io_analog[10] vssa1 6.83fF
C30 io_analog[9] vssa1 6.83fF
C31 m4_204098_586508# vssa1 67.88fF **FLOATING
C32 m4_186716_584374# vssa1 63.83fF **FLOATING
C33 m3_417434_589490# vssa1 3.42fF **FLOATING
C34 io_analog[2] vssa1 20.77fF
C35 L2 vssa1 104.13fF
C36 io_analog[3] vssa1 20.99fF
C37 L1 vssa1 110.57fF
C38 compaartor_v4_0/latch_2_0/inv_W2_1/Vin vssa1 2.76fF
C39 compaartor_v4_0/latch_2_0/inv_W2_0/Vin vssa1 3.67fF
C40 compaartor_v4_0/m1_n58_544# vssa1 2.02fF
C41 io_analog[5] vssa1 339.85fF
C42 io_analog[6] vssa1 358.66fF
C43 compaartor_v4_0/Outp vssa1 111.06fF
C44 compaartor_v4_0/Outn vssa1 104.23fF
C45 CB vssa1 3.33fF
C46 io_analog[7] vssa1 355.98fF
C47 compaartor_v4_0/CLK vssa1 17.42fF
C48 vccd1 vssa1 1929.80fF
C49 io_analog[8] vssa1 383.53fF
.ends

